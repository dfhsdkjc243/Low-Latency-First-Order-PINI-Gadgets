module AESSbox_PINI(
input clk,
input [7:0] sbin0,
input [7:0] sbin1,
input [133:0] ran,
output [7:0] sbout0,
output [7:0] sbout1
);



// wire [7:0] at0_out0,at0_out1,sb0_out0,sb0_out1,at1_out0,at1_out1;



// AffineTrans0_PINI at0(
// .clk(clk),
// .ATin0(a0b0c0d0e0f0g0h0),
// .ATin1(a1b1c1d1e1f1g1h1),
// .ATout0(at0_out0),
// .ATout1(at0_out1)

// );

// TestSbox_trivialopt_l4_PINI sb0(
// .clk(clk),
// .a0b0c0d0e0f0g0h0(at0_out0),
// .a1b1c1d1e1f1g1h1(at0_out1),
// .ran(ran),
// .x0y0z0t0m0n0p0q0(sb0_out0),
// .x1y1z1t1m1n1p1q1(sb0_out1)

// );


// AffineTrans1_PINI at1(
// .clk(clk),
// .ATin0(sb0_out0),
// .ATin1(sb0_out1),
// .ATout0(at1_out0),
// .ATout1(at1_out1)

// );

// assign x0y0z0t0m0n0p0q0 = at1_out0;
// assign x1y1z1t1m1n1p1q1 = at1_out1;




wire [7:0] ATin0, ATin1, ATout0, ATout1;

assign sbin0 = ATin0;
assign sbin1 = ATin1;

wire [7:0] matrix0[0:7];
assign {matrix0[0], matrix0[1], matrix0[2], matrix0[3], matrix0[4], matrix0[5], matrix0[6], matrix0[7]} = {8'h7C ,8'h94 ,8'hB6 ,8'h2A ,8'hDD ,8'h54 ,8'h3C ,8'h70 };
wire [7:0] constant0;
assign constant0 = 8'h00 ;



assign ATout0[7:7] = (matrix0[0][7:7]&ATin0[7:7]) ^ (matrix0[0][6:6]&ATin0[6:6]) ^ (matrix0[0][5:5]&ATin0[5:5]) ^ (matrix0[0][4:4]&ATin0[4:4]) ^ (matrix0[0][3:3]&ATin0[3:3]) ^ (matrix0[0][2:2]&ATin0[2:2]) ^ (matrix0[0][1:1]&ATin0[1:1]) ^ (matrix0[0][0:0]&ATin0[0:0]) ^ constant0[7:7]; 
assign ATout0[6:6] = (matrix0[1][7:7]&ATin0[7:7]) ^ (matrix0[1][6:6]&ATin0[6:6]) ^ (matrix0[1][5:5]&ATin0[5:5]) ^ (matrix0[1][4:4]&ATin0[4:4]) ^ (matrix0[1][3:3]&ATin0[3:3]) ^ (matrix0[1][2:2]&ATin0[2:2]) ^ (matrix0[1][1:1]&ATin0[1:1]) ^ (matrix0[1][0:0]&ATin0[0:0]) ^ constant0[6:6]; 
assign ATout0[5:5] = (matrix0[2][7:7]&ATin0[7:7]) ^ (matrix0[2][6:6]&ATin0[6:6]) ^ (matrix0[2][5:5]&ATin0[5:5]) ^ (matrix0[2][4:4]&ATin0[4:4]) ^ (matrix0[2][3:3]&ATin0[3:3]) ^ (matrix0[2][2:2]&ATin0[2:2]) ^ (matrix0[2][1:1]&ATin0[1:1]) ^ (matrix0[2][0:0]&ATin0[0:0]) ^ constant0[5:5]; 
assign ATout0[4:4] = (matrix0[3][7:7]&ATin0[7:7]) ^ (matrix0[3][6:6]&ATin0[6:6]) ^ (matrix0[3][5:5]&ATin0[5:5]) ^ (matrix0[3][4:4]&ATin0[4:4]) ^ (matrix0[3][3:3]&ATin0[3:3]) ^ (matrix0[3][2:2]&ATin0[2:2]) ^ (matrix0[3][1:1]&ATin0[1:1]) ^ (matrix0[3][0:0]&ATin0[0:0]) ^ constant0[4:4]; 
assign ATout0[3:3] = (matrix0[4][7:7]&ATin0[7:7]) ^ (matrix0[4][6:6]&ATin0[6:6]) ^ (matrix0[4][5:5]&ATin0[5:5]) ^ (matrix0[4][4:4]&ATin0[4:4]) ^ (matrix0[4][3:3]&ATin0[3:3]) ^ (matrix0[4][2:2]&ATin0[2:2]) ^ (matrix0[4][1:1]&ATin0[1:1]) ^ (matrix0[4][0:0]&ATin0[0:0]) ^ constant0[3:3]; 
assign ATout0[2:2] = (matrix0[5][7:7]&ATin0[7:7]) ^ (matrix0[5][6:6]&ATin0[6:6]) ^ (matrix0[5][5:5]&ATin0[5:5]) ^ (matrix0[5][4:4]&ATin0[4:4]) ^ (matrix0[5][3:3]&ATin0[3:3]) ^ (matrix0[5][2:2]&ATin0[2:2]) ^ (matrix0[5][1:1]&ATin0[1:1]) ^ (matrix0[5][0:0]&ATin0[0:0]) ^ constant0[2:2]; 
assign ATout0[1:1] = (matrix0[6][7:7]&ATin0[7:7]) ^ (matrix0[6][6:6]&ATin0[6:6]) ^ (matrix0[6][5:5]&ATin0[5:5]) ^ (matrix0[6][4:4]&ATin0[4:4]) ^ (matrix0[6][3:3]&ATin0[3:3]) ^ (matrix0[6][2:2]&ATin0[2:2]) ^ (matrix0[6][1:1]&ATin0[1:1]) ^ (matrix0[6][0:0]&ATin0[0:0]) ^ constant0[1:1]; 
assign ATout0[0:0] = (matrix0[7][7:7]&ATin0[7:7]) ^ (matrix0[7][6:6]&ATin0[6:6]) ^ (matrix0[7][5:5]&ATin0[5:5]) ^ (matrix0[7][4:4]&ATin0[4:4]) ^ (matrix0[7][3:3]&ATin0[3:3]) ^ (matrix0[7][2:2]&ATin0[2:2]) ^ (matrix0[7][1:1]&ATin0[1:1]) ^ (matrix0[7][0:0]&ATin0[0:0]) ^ constant0[0:0]; 


assign ATout1[7:7] = (matrix0[0][7:7]&ATin1[7:7]) ^ (matrix0[0][6:6]&ATin1[6:6]) ^ (matrix0[0][5:5]&ATin1[5:5]) ^ (matrix0[0][4:4]&ATin1[4:4]) ^ (matrix0[0][3:3]&ATin1[3:3]) ^ (matrix0[0][2:2]&ATin1[2:2]) ^ (matrix0[0][1:1]&ATin1[1:1]) ^ (matrix0[0][0:0]&ATin1[0:0]); 
assign ATout1[6:6] = (matrix0[1][7:7]&ATin1[7:7]) ^ (matrix0[1][6:6]&ATin1[6:6]) ^ (matrix0[1][5:5]&ATin1[5:5]) ^ (matrix0[1][4:4]&ATin1[4:4]) ^ (matrix0[1][3:3]&ATin1[3:3]) ^ (matrix0[1][2:2]&ATin1[2:2]) ^ (matrix0[1][1:1]&ATin1[1:1]) ^ (matrix0[1][0:0]&ATin1[0:0]); 
assign ATout1[5:5] = (matrix0[2][7:7]&ATin1[7:7]) ^ (matrix0[2][6:6]&ATin1[6:6]) ^ (matrix0[2][5:5]&ATin1[5:5]) ^ (matrix0[2][4:4]&ATin1[4:4]) ^ (matrix0[2][3:3]&ATin1[3:3]) ^ (matrix0[2][2:2]&ATin1[2:2]) ^ (matrix0[2][1:1]&ATin1[1:1]) ^ (matrix0[2][0:0]&ATin1[0:0]); 
assign ATout1[4:4] = (matrix0[3][7:7]&ATin1[7:7]) ^ (matrix0[3][6:6]&ATin1[6:6]) ^ (matrix0[3][5:5]&ATin1[5:5]) ^ (matrix0[3][4:4]&ATin1[4:4]) ^ (matrix0[3][3:3]&ATin1[3:3]) ^ (matrix0[3][2:2]&ATin1[2:2]) ^ (matrix0[3][1:1]&ATin1[1:1]) ^ (matrix0[3][0:0]&ATin1[0:0]); 
assign ATout1[3:3] = (matrix0[4][7:7]&ATin1[7:7]) ^ (matrix0[4][6:6]&ATin1[6:6]) ^ (matrix0[4][5:5]&ATin1[5:5]) ^ (matrix0[4][4:4]&ATin1[4:4]) ^ (matrix0[4][3:3]&ATin1[3:3]) ^ (matrix0[4][2:2]&ATin1[2:2]) ^ (matrix0[4][1:1]&ATin1[1:1]) ^ (matrix0[4][0:0]&ATin1[0:0]); 
assign ATout1[2:2] = (matrix0[5][7:7]&ATin1[7:7]) ^ (matrix0[5][6:6]&ATin1[6:6]) ^ (matrix0[5][5:5]&ATin1[5:5]) ^ (matrix0[5][4:4]&ATin1[4:4]) ^ (matrix0[5][3:3]&ATin1[3:3]) ^ (matrix0[5][2:2]&ATin1[2:2]) ^ (matrix0[5][1:1]&ATin1[1:1]) ^ (matrix0[5][0:0]&ATin1[0:0]); 
assign ATout1[1:1] = (matrix0[6][7:7]&ATin1[7:7]) ^ (matrix0[6][6:6]&ATin1[6:6]) ^ (matrix0[6][5:5]&ATin1[5:5]) ^ (matrix0[6][4:4]&ATin1[4:4]) ^ (matrix0[6][3:3]&ATin1[3:3]) ^ (matrix0[6][2:2]&ATin1[2:2]) ^ (matrix0[6][1:1]&ATin1[1:1]) ^ (matrix0[6][0:0]&ATin1[0:0]); 
assign ATout1[0:0] = (matrix0[7][7:7]&ATin1[7:7]) ^ (matrix0[7][6:6]&ATin1[6:6]) ^ (matrix0[7][5:5]&ATin1[5:5]) ^ (matrix0[7][4:4]&ATin1[4:4]) ^ (matrix0[7][3:3]&ATin1[3:3]) ^ (matrix0[7][2:2]&ATin1[2:2]) ^ (matrix0[7][1:1]&ATin1[1:1]) ^ (matrix0[7][0:0]&ATin1[0:0]); 



wire [7:0] a0b0c0d0e0f0g0h0, a1b1c1d1e1f1g1h1, x0y0z0t0m0n0p0q0, x1y1z1t1m1n1p1q1;


assign a0b0c0d0e0f0g0h0 = ATout0;
assign a1b1c1d1e1f1g1h1 = ATout1;

wire a0,b0,c0,d0,e0,f0,g0,h0;
wire a1,b1,c1,d1,e1,f1,g1,h1;
wire r0m, r1m, r2m, r3m, r4m, r5m, r6m, r7m, r8m, r9m, r10m, r11m, r12m, r13m, r14m, r15m, r16m, r17m, r18m, r19m, r20m, r21m, r22m, r23m, r24m, r25m, r26m, r27m, r28m, r29m, r30m, r31m, r32m, r33m, r34m, r35m, r36m, r37m, r38m, r39m, r40m, r41m, r42m, r43m, r44m, r45m, r46m, r47m, r48m, r49m, r50m, r51m, r52m, r53m, r54m, r55m, r56m, r57m, r58m, r59m, r60m, r61m, r62m, r63m, r64m, r65m, r66m, r67m, r68m, r69m, r70m, r71m, r72m, r73m, r74m, r75m, r76m, r77m, r78m, r79m, r80m, r81m, r82m, r83m, r84m, r85m, r86m, r87m, r88m, r89m, r90m, r91m, r92m, r93m, r94m, r95m, r96m, r97m, r98m, r99m, r100m, r101m, r102m, r103m, r104m, r105m, r106m, r107m, r108m, r109m, r110m, r111m, r112m, r113m, r114m, r115m, r116m, r117m, r118m, r119m, r120m, r121m, r122m, r123m, r124m, r125m, r126m, r127m, r128m, r129m, r130m, r131m, r132m, r133m;

assign {h0,g0,f0,e0,d0,c0,b0,a0} = a0b0c0d0e0f0g0h0;
assign {h1,g1,f1,e1,d1,c1,b1,a1} = a1b1c1d1e1f1g1h1;
assign {r0m, r1m, r2m, r3m, r4m, r5m, r6m, r7m, r8m, r9m, r10m, r11m, r12m, r13m, r14m, r15m, r16m, r17m, r18m, r19m, r20m, r21m, r22m, r23m, r24m, r25m, r26m, r27m, r28m, r29m, r30m, r31m, r32m, r33m, r34m, r35m, r36m, r37m, r38m, r39m, r40m, r41m, r42m, r43m, r44m, r45m, r46m, r47m, r48m, r49m, r50m, r51m, r52m, r53m, r54m, r55m, r56m, r57m, r58m, r59m, r60m, r61m, r62m, r63m, r64m, r65m, r66m, r67m, r68m, r69m, r70m, r71m, r72m, r73m, r74m, r75m, r76m, r77m, r78m, r79m, r80m, r81m, r82m, r83m, r84m, r85m, r86m, r87m, r88m, r89m, r90m, r91m, r92m, r93m, r94m, r95m, r96m, r97m, r98m, r99m, r100m, r101m, r102m, r103m, r104m, r105m, r106m, r107m, r108m, r109m, r110m, r111m, r112m, r113m, r114m, r115m, r116m, r117m, r118m, r119m, r120m, r121m, r122m, r123m, r124m, r125m, r126m, r127m, r128m, r129m, r130m, r131m, r132m, r133m} = ran;

reg reg_0_0, reg_0_1, reg_0_2, reg_0_3, reg_0_4, reg_0_5, reg_0_6, reg_0_7, reg_0_8, reg_0_9, reg_0_10, reg_0_11, reg_0_12, reg_0_13, reg_0_14, reg_0_15, reg_0_16, reg_0_17, reg_0_18, reg_0_19, reg_0_20, reg_0_21, reg_0_22, reg_0_23, reg_0_24, reg_0_25, reg_0_26, reg_0_27, reg_0_28, reg_0_29, reg_0_30, reg_0_31, reg_0_32, reg_0_33, reg_0_34, reg_0_35, reg_0_36, reg_0_37, reg_0_38, reg_0_39, reg_0_40, reg_0_41, reg_0_42, reg_0_43, reg_0_44, reg_0_45, reg_0_46, reg_0_47, reg_0_48, reg_0_49, reg_0_50, reg_0_51, reg_0_52, reg_0_53, reg_0_54, reg_0_55, reg_0_56, reg_0_57, reg_0_58, reg_0_59, reg_0_60, reg_0_61, reg_0_62, reg_0_63, reg_0_64, reg_0_65, reg_0_66, reg_0_67, reg_0_68, reg_0_69, reg_0_70, reg_0_71, reg_0_72, reg_0_73, reg_0_74, reg_0_75, reg_0_76, reg_0_77, reg_0_78, reg_0_79, reg_0_80, reg_0_81, reg_0_82, reg_0_83, reg_0_84, reg_0_85, reg_0_86, reg_0_87, reg_0_88, reg_0_89, reg_0_90, reg_0_91, reg_0_92, reg_0_93, reg_0_94, reg_0_95, reg_0_96, reg_0_97, reg_0_98, reg_0_99, reg_0_100, reg_0_101, reg_0_102, reg_0_103, reg_0_104, reg_0_105, reg_0_106, reg_0_107, reg_0_108, reg_0_109, reg_0_110, reg_0_111, reg_0_112, reg_0_113, reg_0_114, reg_0_115, reg_0_116, reg_0_117, reg_0_118, reg_0_119, reg_0_120, reg_0_121, reg_0_122, reg_0_123, reg_0_124, reg_0_125, reg_0_126, reg_0_127, reg_0_128, reg_0_129, reg_0_130, reg_0_131, reg_0_132, reg_0_133, reg_0_134, reg_0_135, reg_0_136, reg_0_137, reg_0_138, reg_0_139, reg_0_140, reg_0_141;
reg reg_1_0, reg_1_1, reg_1_2, reg_1_3, reg_1_4, reg_1_5, reg_1_6, reg_1_7, reg_1_8, reg_1_9, reg_1_10, reg_1_11, reg_1_12, reg_1_13, reg_1_14, reg_1_15, reg_1_16, reg_1_17, reg_1_18, reg_1_19, reg_1_20, reg_1_21, reg_1_22, reg_1_23, reg_1_24, reg_1_25, reg_1_26, reg_1_27, reg_1_28, reg_1_29, reg_1_30, reg_1_31, reg_1_32, reg_1_33, reg_1_34, reg_1_35, reg_1_36, reg_1_37, reg_1_38, reg_1_39, reg_1_40, reg_1_41, reg_1_42, reg_1_43, reg_1_44, reg_1_45, reg_1_46, reg_1_47, reg_1_48, reg_1_49, reg_1_50, reg_1_51, reg_1_52, reg_1_53, reg_1_54, reg_1_55, reg_1_56, reg_1_57, reg_1_58, reg_1_59, reg_1_60, reg_1_61, reg_1_62, reg_1_63, reg_1_64, reg_1_65, reg_1_66, reg_1_67, reg_1_68, reg_1_69, reg_1_70, reg_1_71, reg_1_72, reg_1_73, reg_1_74, reg_1_75, reg_1_76, reg_1_77, reg_1_78, reg_1_79, reg_1_80, reg_1_81, reg_1_82, reg_1_83, reg_1_84, reg_1_85, reg_1_86, reg_1_87, reg_1_88, reg_1_89, reg_1_90, reg_1_91, reg_1_92, reg_1_93, reg_1_94, reg_1_95, reg_1_96, reg_1_97, reg_1_98, reg_1_99, reg_1_100, reg_1_101, reg_1_102, reg_1_103, reg_1_104, reg_1_105, reg_1_106, reg_1_107, reg_1_108, reg_1_109, reg_1_110, reg_1_111, reg_1_112, reg_1_113, reg_1_114, reg_1_115, reg_1_116, reg_1_117, reg_1_118, reg_1_119, reg_1_120, reg_1_121, reg_1_122, reg_1_123, reg_1_124, reg_1_125, reg_1_126, reg_1_127, reg_1_128, reg_1_129, reg_1_130, reg_1_131, reg_1_132, reg_1_133, reg_1_134, reg_1_135, reg_1_136, reg_1_137, reg_1_138, reg_1_139, reg_1_140, reg_1_141;




wire cdxi0m = (b1 ^ r0m);
wire cdxi1m = (c1 ^ r1m);
wire cdxi2m = (d1 ^ r2m);
wire cdxi3m = (e1 ^ r3m);
wire cdxi4m = (f1 ^ r4m);
wire cdxi5m = (g1 ^ r5m);
wire cdxi6m = (h1 ^ r6m);
wire cdxi7m = b1&c1 ^ r7m;
wire cdxi8m = b1&d1 ^ r8m;
wire cdxi9m = b1&e1 ^ r9m;
wire cdxi10m = b1&f1 ^ r10m;
wire cdxi11m = b1&g1 ^ r11m;
wire cdxi12m = b1&h1 ^ r12m;
wire cdxi13m = c1&d1 ^ r13m;
wire cdxi14m = c1&e1 ^ r14m;
wire cdxi15m = c1&f1 ^ r15m;
wire cdxi16m = c1&g1 ^ r16m;
wire cdxi17m = c1&h1 ^ r17m;
wire cdxi18m = d1&e1 ^ r18m;
wire cdxi19m = d1&f1 ^ r19m;
wire cdxi20m = d1&g1 ^ r20m;
wire cdxi21m = d1&h1 ^ r21m;
wire cdxi22m = e1&f1 ^ r22m;
wire cdxi23m = e1&g1 ^ r23m;
wire cdxi24m = e1&h1 ^ r24m;
wire cdxi25m = f1&g1 ^ r25m;
wire cdxi26m = f1&h1 ^ r26m;
wire cdxi27m = g1&h1 ^ r27m;
wire cdxi28m = b1&c1&d1 ^ r28m;
wire cdxi29m = b1&c1&e1 ^ r29m;
wire cdxi30m = b1&c1&f1 ^ r30m;
wire cdxi31m = b1&c1&g1 ^ r31m;
wire cdxi32m = b1&c1&h1 ^ r32m;
wire cdxi33m = b1&d1&e1 ^ r33m;
wire cdxi34m = b1&d1&f1 ^ r34m;
wire cdxi35m = b1&d1&g1 ^ r35m;
wire cdxi36m = b1&d1&h1 ^ r36m;
wire cdxi37m = b1&e1&f1 ^ r37m;
wire cdxi38m = b1&e1&g1 ^ r38m;
wire cdxi39m = b1&e1&h1 ^ r39m;
wire cdxi40m = b1&f1&g1 ^ r40m;
wire cdxi41m = b1&f1&h1 ^ r41m;
wire cdxi42m = b1&g1&h1 ^ r42m;
wire cdxi43m = c1&d1&e1 ^ r43m;
wire cdxi44m = c1&d1&f1 ^ r44m;
wire cdxi45m = c1&d1&g1 ^ r45m;
wire cdxi46m = c1&d1&h1 ^ r46m;
wire cdxi47m = c1&e1&f1 ^ r47m;
wire cdxi48m = c1&e1&g1 ^ r48m;
wire cdxi49m = c1&e1&h1 ^ r49m;
wire cdxi50m = c1&f1&g1 ^ r50m;
wire cdxi51m = c1&f1&h1 ^ r51m;
wire cdxi52m = c1&g1&h1 ^ r52m;
wire cdxi53m = d1&e1&f1 ^ r53m;
wire cdxi54m = d1&e1&g1 ^ r54m;
wire cdxi55m = d1&e1&h1 ^ r55m;
wire cdxi56m = d1&f1&g1 ^ r56m;
wire cdxi57m = d1&f1&h1 ^ r57m;
wire cdxi58m = d1&g1&h1 ^ r58m;
wire cdxi59m = e1&f1&g1 ^ r59m;
wire cdxi60m = e1&f1&h1 ^ r60m;
wire cdxi61m = e1&g1&h1 ^ r61m;
wire cdxi62m = f1&g1&h1 ^ r62m;
wire cdxi63m = b1&c1&d1&e1 ^ r63m;
wire cdxi64m = b1&c1&d1&f1 ^ r64m;
wire cdxi65m = b1&c1&d1&g1 ^ r65m;
wire cdxi66m = b1&c1&d1&h1 ^ r66m;
wire cdxi67m = b1&c1&e1&f1 ^ r67m;
wire cdxi68m = b1&c1&e1&g1 ^ r68m;
wire cdxi69m = b1&c1&e1&h1 ^ r69m;
wire cdxi70m = b1&c1&f1&g1 ^ r70m;
wire cdxi71m = b1&c1&f1&h1 ^ r71m;
wire cdxi72m = b1&c1&g1&h1 ^ r72m;
wire cdxi73m = b1&d1&e1&f1 ^ r73m;
wire cdxi74m = b1&d1&e1&g1 ^ r74m;
wire cdxi75m = b1&d1&e1&h1 ^ r75m;
wire cdxi76m = b1&d1&f1&g1 ^ r76m;
wire cdxi77m = b1&d1&f1&h1 ^ r77m;
wire cdxi78m = b1&d1&g1&h1 ^ r78m;
wire cdxi79m = b1&e1&f1&g1 ^ r79m;
wire cdxi80m = b1&e1&f1&h1 ^ r80m;
wire cdxi81m = b1&e1&g1&h1 ^ r81m;
wire cdxi82m = b1&f1&g1&h1 ^ r82m;
wire cdxi83m = c1&d1&e1&f1 ^ r83m;
wire cdxi84m = c1&d1&e1&g1 ^ r84m;
wire cdxi85m = c1&d1&e1&h1 ^ r85m;
wire cdxi86m = c1&d1&f1&g1 ^ r86m;
wire cdxi87m = c1&d1&f1&h1 ^ r87m;
wire cdxi88m = c1&d1&g1&h1 ^ r88m;
wire cdxi89m = c1&e1&f1&g1 ^ r89m;
wire cdxi90m = c1&e1&f1&h1 ^ r90m;
wire cdxi91m = c1&e1&g1&h1 ^ r91m;
wire cdxi92m = c1&f1&g1&h1 ^ r92m;
wire cdxi93m = d1&e1&f1&g1 ^ r93m;
wire cdxi94m = d1&e1&f1&h1 ^ r94m;
wire cdxi95m = d1&e1&g1&h1 ^ r95m;
wire cdxi96m = d1&f1&g1&h1 ^ r96m;
wire cdxi97m = e1&f1&g1&h1 ^ r97m;
wire cdxi98m = b1&c1&d1&e1&f1 ^ r98m;
wire cdxi99m = b1&c1&d1&e1&g1 ^ r99m;
wire cdxi100m = b1&c1&d1&e1&h1 ^ r100m;
wire cdxi101m = b1&c1&d1&f1&g1 ^ r101m;
wire cdxi102m = b1&c1&d1&f1&h1 ^ r102m;
wire cdxi103m = b1&c1&d1&g1&h1 ^ r103m;
wire cdxi104m = b1&c1&e1&f1&g1 ^ r104m;
wire cdxi105m = b1&c1&e1&f1&h1 ^ r105m;
wire cdxi106m = b1&c1&e1&g1&h1 ^ r106m;
wire cdxi107m = b1&c1&f1&g1&h1 ^ r107m;
wire cdxi108m = b1&d1&e1&f1&g1 ^ r108m;
wire cdxi109m = b1&d1&e1&f1&h1 ^ r109m;
wire cdxi110m = b1&d1&e1&g1&h1 ^ r110m;
wire cdxi111m = b1&d1&f1&g1&h1 ^ r111m;
wire cdxi112m = b1&e1&f1&g1&h1 ^ r112m;
wire cdxi113m = c1&d1&e1&f1&g1 ^ r113m;
wire cdxi114m = c1&d1&e1&f1&h1 ^ r114m;
wire cdxi115m = c1&d1&e1&g1&h1 ^ r115m;
wire cdxi116m = c1&d1&f1&g1&h1 ^ r116m;
wire cdxi117m = c1&e1&f1&g1&h1 ^ r117m;
wire cdxi118m = d1&e1&f1&g1&h1 ^ r118m;
wire cdxi119m = b1&c1&d1&e1&f1&g1 ^ r119m;
wire cdxi120m = b1&c1&d1&e1&f1&h1 ^ r120m;
wire cdxi121m = b1&c1&d1&e1&g1&h1 ^ r121m;
wire cdxi122m = b1&c1&d1&f1&g1&h1 ^ r122m;
wire cdxi123m = b1&c1&e1&f1&g1&h1 ^ r123m;
wire cdxi124m = b1&d1&e1&f1&g1&h1 ^ r124m;
wire cdxi125m = c1&d1&e1&f1&g1&h1 ^ r125m;
wire cdxi126m = 1&1 ^ a0 ^ b0 ^ c0 ^ f0;
wire cdxi127m = b0 ^ r0m;
wire cdxi128m = (cdxi127m);
wire cdxi129m = a0&cdxi128m;
wire cdxi130m = (reg_0_8);
wire cdxi131m = (cdxi130m);
wire cdxi132m = reg_0_0&cdxi131m;
wire cdxi133m = c0 ^ r1m;
wire cdxi134m = (cdxi133m);
wire cdxi135m = a0&cdxi134m;
wire cdxi136m = (reg_0_9);
wire cdxi137m = (cdxi136m);
wire cdxi138m = reg_0_0&cdxi137m;
wire cdxi139m = d0 ^ r2m;
wire cdxi140m = (cdxi139m);
wire cdxi141m = a0&cdxi140m;
wire cdxi142m = (reg_0_10);
wire cdxi143m = (cdxi142m);
wire cdxi144m = reg_0_0&cdxi143m;
wire cdxi145m = e0 ^ r3m;
wire cdxi146m = (cdxi145m);
wire cdxi147m = a0&cdxi146m;
wire cdxi148m = (reg_0_11);
wire cdxi149m = (cdxi148m);
wire cdxi150m = reg_0_0&cdxi149m;
wire cdxi151m = f0 ^ r4m;
wire cdxi152m = (cdxi151m);
wire cdxi153m = a0&cdxi152m;
wire cdxi154m = (reg_0_12);
wire cdxi155m = (cdxi154m);
wire cdxi156m = reg_0_0&cdxi155m;
wire cdxi157m = g0 ^ r5m;
wire cdxi158m = (cdxi157m);
wire cdxi159m = a0&cdxi158m;
wire cdxi160m = (reg_0_13);
wire cdxi161m = (cdxi160m);
wire cdxi162m = reg_0_0&cdxi161m;
wire cdxi163m = b0&cdxi140m;
wire cdxi164m = reg_0_1&cdxi143m;
wire cdxi165m = b0&cdxi158m;
wire cdxi166m = reg_0_1&cdxi161m;
wire cdxi167m = h0 ^ r6m;
wire cdxi168m = (cdxi167m);
wire cdxi169m = b0&cdxi168m;
wire cdxi170m = (reg_0_14);
wire cdxi171m = (cdxi170m);
wire cdxi172m = reg_0_1&cdxi171m;
wire cdxi173m = c0&cdxi158m;
wire cdxi174m = reg_0_2&cdxi161m;
wire cdxi175m = d0&cdxi152m;
wire cdxi176m = reg_0_3&cdxi155m;
wire cdxi177m = e0&cdxi158m;
wire cdxi178m = reg_0_4&cdxi161m;
wire cdxi179m = e0&cdxi168m;
wire cdxi180m = reg_0_4&cdxi171m;
wire cdxi181m = f0&cdxi158m;
wire cdxi182m = reg_0_5&cdxi161m;
wire cdxi183m = b0&d0 ^ r8m;
wire cdxi184m = d0;
wire cdxi185m = b0;
wire cdxi186m = cdxi184m&r0m;
wire cdxi187m = cdxi185m&r2m;
wire cdxi188m = (cdxi183m ^ cdxi186m ^ cdxi187m);
wire cdxi189m = a0&cdxi188m;
wire cdxi190m = (reg_0_16);
wire cdxi191m = reg_0_3&cdxi130m;
wire cdxi192m = reg_0_1&cdxi142m;
wire cdxi193m = (cdxi191m ^ cdxi192m ^ cdxi190m);
wire cdxi194m = reg_0_0&cdxi193m;
wire cdxi195m = cdxi185m&e0 ^ r9m;
wire cdxi196m = e0;
wire cdxi197m = cdxi196m&r0m;
wire cdxi198m = cdxi185m&r3m;
wire cdxi199m = (cdxi195m ^ cdxi197m ^ cdxi198m);
wire cdxi200m = a0&cdxi199m;
wire cdxi201m = (reg_0_17);
wire cdxi202m = reg_0_4&cdxi130m;
wire cdxi203m = reg_0_1&cdxi148m;
wire cdxi204m = (cdxi202m ^ cdxi203m ^ cdxi201m);
wire cdxi205m = reg_0_0&cdxi204m;
wire cdxi206m = cdxi185m&h0 ^ r12m;
wire cdxi207m = h0;
wire cdxi208m = cdxi207m&r0m;
wire cdxi209m = cdxi185m&r6m;
wire cdxi210m = (cdxi206m ^ cdxi208m ^ cdxi209m);
wire cdxi211m = a0&cdxi210m;
wire cdxi212m = (reg_0_20);
wire cdxi213m = reg_0_7&cdxi130m;
wire cdxi214m = reg_0_1&cdxi170m;
wire cdxi215m = (cdxi213m ^ cdxi214m ^ cdxi212m);
wire cdxi216m = reg_0_0&cdxi215m;
wire cdxi217m = c0&g0 ^ r16m;
wire cdxi218m = g0;
wire cdxi219m = c0;
wire cdxi220m = cdxi218m&r1m;
wire cdxi221m = cdxi219m&r5m;
wire cdxi222m = (cdxi217m ^ cdxi220m ^ cdxi221m);
wire cdxi223m = a0&cdxi222m;
wire cdxi224m = (reg_0_24);
wire cdxi225m = reg_0_6&cdxi136m;
wire cdxi226m = reg_0_2&cdxi160m;
wire cdxi227m = (cdxi225m ^ cdxi226m ^ cdxi224m);
wire cdxi228m = reg_0_0&cdxi227m;
wire cdxi229m = cdxi184m&cdxi207m ^ r21m;
wire cdxi230m = cdxi207m&r2m;
wire cdxi231m = cdxi184m&r6m;
wire cdxi232m = (cdxi229m ^ cdxi230m ^ cdxi231m);
wire cdxi233m = a0&cdxi232m;
wire cdxi234m = (reg_0_29);
wire cdxi235m = reg_0_7&cdxi142m;
wire cdxi236m = reg_0_3&cdxi170m;
wire cdxi237m = (cdxi235m ^ cdxi236m ^ cdxi234m);
wire cdxi238m = reg_0_0&cdxi237m;
wire cdxi239m = cdxi196m&f0 ^ r22m;
wire cdxi240m = f0;
wire cdxi241m = cdxi240m&r3m;
wire cdxi242m = cdxi196m&r4m;
wire cdxi243m = (cdxi239m ^ cdxi241m ^ cdxi242m);
wire cdxi244m = a0&cdxi243m;
wire cdxi245m = (reg_0_30);
wire cdxi246m = reg_0_5&cdxi148m;
wire cdxi247m = reg_0_4&cdxi154m;
wire cdxi248m = (cdxi246m ^ cdxi247m ^ cdxi245m);
wire cdxi249m = reg_0_0&cdxi248m;
wire cdxi250m = cdxi240m&cdxi218m ^ r25m;
wire cdxi251m = cdxi218m&r4m;
wire cdxi252m = cdxi240m&r5m;
wire cdxi253m = (cdxi250m ^ cdxi251m ^ cdxi252m);
wire cdxi254m = a0&cdxi253m;
wire cdxi255m = (reg_0_33);
wire cdxi256m = reg_0_6&cdxi154m;
wire cdxi257m = reg_0_5&cdxi160m;
wire cdxi258m = (cdxi256m ^ cdxi257m ^ cdxi255m);
wire cdxi259m = reg_0_0&cdxi258m;
wire cdxi260m = cdxi240m&cdxi207m ^ r26m;
wire cdxi261m = cdxi207m&r4m;
wire cdxi262m = cdxi240m&r6m;
wire cdxi263m = (cdxi260m ^ cdxi261m ^ cdxi262m);
wire cdxi264m = a0&cdxi263m;
wire cdxi265m = (reg_0_34);
wire cdxi266m = reg_0_7&cdxi154m;
wire cdxi267m = reg_0_5&cdxi170m;
wire cdxi268m = (cdxi266m ^ cdxi267m ^ cdxi265m);
wire cdxi269m = reg_0_0&cdxi268m;
wire cdxi270m = cdxi219m&cdxi207m ^ r17m;
wire cdxi271m = cdxi207m&r1m;
wire cdxi272m = cdxi219m&r6m;
wire cdxi273m = (cdxi270m ^ cdxi271m ^ cdxi272m);
wire cdxi274m = cdxi185m&cdxi273m;
wire cdxi275m = (reg_0_25);
wire cdxi276m = reg_0_7&cdxi136m;
wire cdxi277m = reg_0_2&cdxi170m;
wire cdxi278m = (cdxi276m ^ cdxi277m ^ cdxi275m);
wire cdxi279m = reg_0_1&cdxi278m;
wire cdxi280m = cdxi184m&cdxi196m ^ r18m;
wire cdxi281m = cdxi196m&r2m;
wire cdxi282m = cdxi184m&r3m;
wire cdxi283m = (cdxi280m ^ cdxi281m ^ cdxi282m);
wire cdxi284m = cdxi185m&cdxi283m;
wire cdxi285m = (reg_0_26);
wire cdxi286m = reg_0_4&cdxi142m;
wire cdxi287m = reg_0_3&cdxi148m;
wire cdxi288m = (cdxi286m ^ cdxi287m ^ cdxi285m);
wire cdxi289m = reg_0_1&cdxi288m;
wire cdxi290m = cdxi184m&cdxi218m ^ r20m;
wire cdxi291m = cdxi218m&r2m;
wire cdxi292m = cdxi184m&r5m;
wire cdxi293m = (cdxi290m ^ cdxi291m ^ cdxi292m);
wire cdxi294m = cdxi185m&cdxi293m;
wire cdxi295m = (reg_0_28);
wire cdxi296m = reg_0_6&cdxi142m;
wire cdxi297m = reg_0_3&cdxi160m;
wire cdxi298m = (cdxi296m ^ cdxi297m ^ cdxi295m);
wire cdxi299m = reg_0_1&cdxi298m;
wire cdxi300m = cdxi196m&cdxi218m ^ r23m;
wire cdxi301m = cdxi218m&r3m;
wire cdxi302m = cdxi196m&r5m;
wire cdxi303m = (cdxi300m ^ cdxi301m ^ cdxi302m);
wire cdxi304m = cdxi185m&cdxi303m;
wire cdxi305m = (reg_0_31);
wire cdxi306m = reg_0_6&cdxi148m;
wire cdxi307m = reg_0_4&cdxi160m;
wire cdxi308m = (cdxi306m ^ cdxi307m ^ cdxi305m);
wire cdxi309m = reg_0_1&cdxi308m;
wire cdxi310m = cdxi184m&cdxi240m ^ r19m;
wire cdxi311m = cdxi240m&r2m;
wire cdxi312m = cdxi184m&r4m;
wire cdxi313m = (cdxi310m ^ cdxi311m ^ cdxi312m);
wire cdxi314m = cdxi219m&cdxi313m;
wire cdxi315m = (reg_0_27);
wire cdxi316m = reg_0_5&cdxi142m;
wire cdxi317m = reg_0_3&cdxi154m;
wire cdxi318m = (cdxi316m ^ cdxi317m ^ cdxi315m);
wire cdxi319m = reg_0_2&cdxi318m;
wire cdxi320m = cdxi219m&cdxi232m;
wire cdxi321m = reg_0_2&cdxi237m;
wire cdxi322m = cdxi219m&cdxi303m;
wire cdxi323m = reg_0_2&cdxi308m;
wire cdxi324m = cdxi196m&cdxi207m ^ r24m;
wire cdxi325m = cdxi207m&r3m;
wire cdxi326m = cdxi196m&r6m;
wire cdxi327m = (cdxi324m ^ cdxi325m ^ cdxi326m);
wire cdxi328m = cdxi219m&cdxi327m;
wire cdxi329m = (reg_0_32);
wire cdxi330m = reg_0_7&cdxi148m;
wire cdxi331m = reg_0_4&cdxi170m;
wire cdxi332m = (cdxi330m ^ cdxi331m ^ cdxi329m);
wire cdxi333m = reg_0_2&cdxi332m;
wire cdxi334m = cdxi219m&cdxi253m;
wire cdxi335m = reg_0_2&cdxi258m;
wire cdxi336m = cdxi218m&cdxi207m ^ r27m;
wire cdxi337m = cdxi207m&r5m;
wire cdxi338m = cdxi218m&r6m;
wire cdxi339m = (cdxi336m ^ cdxi337m ^ cdxi338m);
wire cdxi340m = cdxi219m&cdxi339m;
wire cdxi341m = (reg_0_35);
wire cdxi342m = reg_0_7&cdxi160m;
wire cdxi343m = reg_0_6&cdxi170m;
wire cdxi344m = (cdxi342m ^ cdxi343m ^ cdxi341m);
wire cdxi345m = reg_0_2&cdxi344m;
wire cdxi346m = cdxi184m&cdxi243m;
wire cdxi347m = reg_0_3&cdxi248m;
wire cdxi348m = cdxi184m&cdxi303m;
wire cdxi349m = reg_0_3&cdxi308m;
wire cdxi350m = cdxi184m&cdxi327m;
wire cdxi351m = reg_0_3&cdxi332m;
wire cdxi352m = cdxi184m&cdxi253m;
wire cdxi353m = reg_0_3&cdxi258m;
wire cdxi354m = cdxi184m&cdxi263m;
wire cdxi355m = reg_0_3&cdxi268m;
wire cdxi356m = cdxi196m&cdxi253m;
wire cdxi357m = reg_0_4&cdxi258m;
wire cdxi358m = cdxi196m&cdxi263m;
wire cdxi359m = reg_0_4&cdxi268m;
wire cdxi360m = cdxi185m&cdxi219m&cdxi184m ^ r28m;
wire cdxi361m = cdxi219m&cdxi184m;
wire cdxi362m = cdxi185m&cdxi184m;
wire cdxi363m = cdxi185m&cdxi219m;
wire cdxi364m = cdxi219m&cdxi186m;
wire cdxi365m = cdxi362m&r1m;
wire cdxi366m = cdxi363m&r2m;
wire cdxi367m = cdxi184m&r7m;
wire cdxi368m = cdxi219m&r8m;
wire cdxi369m = cdxi185m&r13m;
wire cdxi370m = (cdxi360m ^ cdxi364m ^ cdxi365m ^ cdxi366m ^ cdxi367m ^ cdxi368m ^ cdxi369m);
wire cdxi371m = a0&cdxi370m;
wire cdxi372m = (reg_0_15);
wire cdxi373m = (reg_0_21);
wire cdxi374m = (reg_0_36);
wire cdxi375m = reg_0_2&cdxi191m;
wire cdxi376m = reg_0_1&reg_0_3&cdxi136m;
wire cdxi377m = reg_0_1&reg_0_2&cdxi142m;
wire cdxi378m = reg_0_3&cdxi372m;
wire cdxi379m = reg_0_2&cdxi190m;
wire cdxi380m = reg_0_1&cdxi373m;
wire cdxi381m = (cdxi375m ^ cdxi376m ^ cdxi377m ^ cdxi378m ^ cdxi379m ^ cdxi380m ^ cdxi374m);
wire cdxi382m = reg_0_0&cdxi381m;
wire cdxi383m = cdxi363m&cdxi218m ^ r31m;
wire cdxi384m = cdxi219m&cdxi218m;
wire cdxi385m = cdxi185m&cdxi218m;
wire cdxi386m = cdxi384m&r0m;
wire cdxi387m = cdxi185m&cdxi220m;
wire cdxi388m = cdxi185m&cdxi221m;
wire cdxi389m = cdxi218m&r7m;
wire cdxi390m = cdxi219m&r11m;
wire cdxi391m = cdxi185m&r16m;
wire cdxi392m = (cdxi383m ^ cdxi386m ^ cdxi387m ^ cdxi388m ^ cdxi389m ^ cdxi390m ^ cdxi391m);
wire cdxi393m = a0&cdxi392m;
wire cdxi394m = (reg_0_19);
wire cdxi395m = (reg_0_39);
wire cdxi396m = reg_0_2&reg_0_6&cdxi130m;
wire cdxi397m = reg_0_1&cdxi225m;
wire cdxi398m = reg_0_1&cdxi226m;
wire cdxi399m = reg_0_6&cdxi372m;
wire cdxi400m = reg_0_2&cdxi394m;
wire cdxi401m = reg_0_1&cdxi224m;
wire cdxi402m = (cdxi396m ^ cdxi397m ^ cdxi398m ^ cdxi399m ^ cdxi400m ^ cdxi401m ^ cdxi395m);
wire cdxi403m = reg_0_0&cdxi402m;
wire cdxi404m = cdxi362m&cdxi196m ^ r33m;
wire cdxi405m = cdxi184m&cdxi196m;
wire cdxi406m = cdxi185m&cdxi196m;
wire cdxi407m = cdxi184m&cdxi197m;
wire cdxi408m = cdxi185m&cdxi281m;
wire cdxi409m = cdxi185m&cdxi282m;
wire cdxi410m = cdxi196m&r8m;
wire cdxi411m = cdxi184m&r9m;
wire cdxi412m = cdxi185m&r18m;
wire cdxi413m = (cdxi404m ^ cdxi407m ^ cdxi408m ^ cdxi409m ^ cdxi410m ^ cdxi411m ^ cdxi412m);
wire cdxi414m = a0&cdxi413m;
wire cdxi415m = (reg_0_41);
wire cdxi416m = reg_0_3&cdxi202m;
wire cdxi417m = reg_0_1&cdxi286m;
wire cdxi418m = reg_0_1&cdxi287m;
wire cdxi419m = reg_0_4&cdxi190m;
wire cdxi420m = reg_0_3&cdxi201m;
wire cdxi421m = reg_0_1&cdxi285m;
wire cdxi422m = (cdxi416m ^ cdxi417m ^ cdxi418m ^ cdxi419m ^ cdxi420m ^ cdxi421m ^ cdxi415m);
wire cdxi423m = reg_0_0&cdxi422m;
wire cdxi424m = cdxi362m&cdxi207m ^ r36m;
wire cdxi425m = cdxi184m&cdxi207m;
wire cdxi426m = cdxi185m&cdxi207m;
wire cdxi427m = cdxi184m&cdxi208m;
wire cdxi428m = cdxi185m&cdxi230m;
wire cdxi429m = cdxi185m&cdxi231m;
wire cdxi430m = cdxi207m&r8m;
wire cdxi431m = cdxi184m&r12m;
wire cdxi432m = cdxi185m&r21m;
wire cdxi433m = (cdxi424m ^ cdxi427m ^ cdxi428m ^ cdxi429m ^ cdxi430m ^ cdxi431m ^ cdxi432m);
wire cdxi434m = a0&cdxi433m;
wire cdxi435m = (reg_0_44);
wire cdxi436m = reg_0_3&cdxi213m;
wire cdxi437m = reg_0_1&cdxi235m;
wire cdxi438m = reg_0_1&cdxi236m;
wire cdxi439m = reg_0_7&cdxi190m;
wire cdxi440m = reg_0_3&cdxi212m;
wire cdxi441m = reg_0_1&cdxi234m;
wire cdxi442m = (cdxi436m ^ cdxi437m ^ cdxi438m ^ cdxi439m ^ cdxi440m ^ cdxi441m ^ cdxi435m);
wire cdxi443m = reg_0_0&cdxi442m;
wire cdxi444m = cdxi406m&cdxi240m ^ r37m;
wire cdxi445m = cdxi196m&cdxi240m;
wire cdxi446m = cdxi185m&cdxi240m;
wire cdxi447m = cdxi445m&r0m;
wire cdxi448m = cdxi185m&cdxi241m;
wire cdxi449m = cdxi185m&cdxi242m;
wire cdxi450m = cdxi240m&r9m;
wire cdxi451m = cdxi196m&r10m;
wire cdxi452m = cdxi185m&r22m;
wire cdxi453m = (cdxi444m ^ cdxi447m ^ cdxi448m ^ cdxi449m ^ cdxi450m ^ cdxi451m ^ cdxi452m);
wire cdxi454m = a0&cdxi453m;
wire cdxi455m = (reg_0_18);
wire cdxi456m = (reg_0_45);
wire cdxi457m = reg_0_4&reg_0_5&cdxi130m;
wire cdxi458m = reg_0_1&cdxi246m;
wire cdxi459m = reg_0_1&cdxi247m;
wire cdxi460m = reg_0_5&cdxi201m;
wire cdxi461m = reg_0_4&cdxi455m;
wire cdxi462m = reg_0_1&cdxi245m;
wire cdxi463m = (cdxi457m ^ cdxi458m ^ cdxi459m ^ cdxi460m ^ cdxi461m ^ cdxi462m ^ cdxi456m);
wire cdxi464m = reg_0_0&cdxi463m;
wire cdxi465m = cdxi406m&cdxi218m ^ r38m;
wire cdxi466m = cdxi196m&cdxi218m;
wire cdxi467m = cdxi466m&r0m;
wire cdxi468m = cdxi185m&cdxi301m;
wire cdxi469m = cdxi185m&cdxi302m;
wire cdxi470m = cdxi218m&r9m;
wire cdxi471m = cdxi196m&r11m;
wire cdxi472m = cdxi185m&r23m;
wire cdxi473m = (cdxi465m ^ cdxi467m ^ cdxi468m ^ cdxi469m ^ cdxi470m ^ cdxi471m ^ cdxi472m);
wire cdxi474m = a0&cdxi473m;
wire cdxi475m = (reg_0_46);
wire cdxi476m = reg_0_4&reg_0_6&cdxi130m;
wire cdxi477m = reg_0_1&cdxi306m;
wire cdxi478m = reg_0_1&cdxi307m;
wire cdxi479m = reg_0_6&cdxi201m;
wire cdxi480m = reg_0_4&cdxi394m;
wire cdxi481m = reg_0_1&cdxi305m;
wire cdxi482m = (cdxi476m ^ cdxi477m ^ cdxi478m ^ cdxi479m ^ cdxi480m ^ cdxi481m ^ cdxi475m);
wire cdxi483m = reg_0_0&cdxi482m;
wire cdxi484m = cdxi446m&cdxi207m ^ r41m;
wire cdxi485m = cdxi240m&cdxi207m;
wire cdxi486m = cdxi240m&cdxi208m;
wire cdxi487m = cdxi185m&cdxi261m;
wire cdxi488m = cdxi185m&cdxi262m;
wire cdxi489m = cdxi207m&r10m;
wire cdxi490m = cdxi240m&r12m;
wire cdxi491m = cdxi185m&r26m;
wire cdxi492m = (cdxi484m ^ cdxi486m ^ cdxi487m ^ cdxi488m ^ cdxi489m ^ cdxi490m ^ cdxi491m);
wire cdxi493m = a0&cdxi492m;
wire cdxi494m = (reg_0_49);
wire cdxi495m = reg_0_5&cdxi213m;
wire cdxi496m = reg_0_1&cdxi266m;
wire cdxi497m = reg_0_1&cdxi267m;
wire cdxi498m = reg_0_7&cdxi455m;
wire cdxi499m = reg_0_5&cdxi212m;
wire cdxi500m = reg_0_1&cdxi265m;
wire cdxi501m = (cdxi495m ^ cdxi496m ^ cdxi497m ^ cdxi498m ^ cdxi499m ^ cdxi500m ^ cdxi494m);
wire cdxi502m = reg_0_0&cdxi501m;
wire cdxi503m = cdxi361m&cdxi196m ^ r43m;
wire cdxi504m = cdxi219m&cdxi196m;
wire cdxi505m = cdxi405m&r1m;
wire cdxi506m = cdxi219m&cdxi281m;
wire cdxi507m = cdxi219m&cdxi282m;
wire cdxi508m = cdxi196m&r13m;
wire cdxi509m = cdxi184m&r14m;
wire cdxi510m = cdxi219m&r18m;
wire cdxi511m = (cdxi503m ^ cdxi505m ^ cdxi506m ^ cdxi507m ^ cdxi508m ^ cdxi509m ^ cdxi510m);
wire cdxi512m = a0&cdxi511m;
wire cdxi513m = (reg_0_22);
wire cdxi514m = (reg_0_51);
wire cdxi515m = reg_0_3&reg_0_4&cdxi136m;
wire cdxi516m = reg_0_2&cdxi286m;
wire cdxi517m = reg_0_2&cdxi287m;
wire cdxi518m = reg_0_4&cdxi373m;
wire cdxi519m = reg_0_3&cdxi513m;
wire cdxi520m = reg_0_2&cdxi285m;
wire cdxi521m = (cdxi515m ^ cdxi516m ^ cdxi517m ^ cdxi518m ^ cdxi519m ^ cdxi520m ^ cdxi514m);
wire cdxi522m = reg_0_0&cdxi521m;
wire cdxi523m = cdxi219m&cdxi445m ^ r47m;
wire cdxi524m = cdxi219m&cdxi240m;
wire cdxi525m = cdxi445m&r1m;
wire cdxi526m = cdxi219m&cdxi241m;
wire cdxi527m = cdxi219m&cdxi242m;
wire cdxi528m = cdxi240m&r14m;
wire cdxi529m = cdxi196m&r15m;
wire cdxi530m = cdxi219m&r22m;
wire cdxi531m = (cdxi523m ^ cdxi525m ^ cdxi526m ^ cdxi527m ^ cdxi528m ^ cdxi529m ^ cdxi530m);
wire cdxi532m = a0&cdxi531m;
wire cdxi533m = (reg_0_23);
wire cdxi534m = (reg_0_55);
wire cdxi535m = reg_0_4&reg_0_5&cdxi136m;
wire cdxi536m = reg_0_2&cdxi246m;
wire cdxi537m = reg_0_2&cdxi247m;
wire cdxi538m = reg_0_5&cdxi513m;
wire cdxi539m = reg_0_4&cdxi533m;
wire cdxi540m = reg_0_2&cdxi245m;
wire cdxi541m = (cdxi535m ^ cdxi536m ^ cdxi537m ^ cdxi538m ^ cdxi539m ^ cdxi540m ^ cdxi534m);
wire cdxi542m = reg_0_0&cdxi541m;
wire cdxi543m = cdxi219m&cdxi466m ^ r48m;
wire cdxi544m = cdxi196m&cdxi220m;
wire cdxi545m = cdxi219m&cdxi301m;
wire cdxi546m = cdxi219m&cdxi302m;
wire cdxi547m = cdxi218m&r14m;
wire cdxi548m = cdxi196m&r16m;
wire cdxi549m = cdxi219m&r23m;
wire cdxi550m = (cdxi543m ^ cdxi544m ^ cdxi545m ^ cdxi546m ^ cdxi547m ^ cdxi548m ^ cdxi549m);
wire cdxi551m = a0&cdxi550m;
wire cdxi552m = (reg_0_56);
wire cdxi553m = reg_0_4&cdxi225m;
wire cdxi554m = reg_0_2&cdxi306m;
wire cdxi555m = reg_0_2&cdxi307m;
wire cdxi556m = reg_0_6&cdxi513m;
wire cdxi557m = reg_0_4&cdxi224m;
wire cdxi558m = reg_0_2&cdxi305m;
wire cdxi559m = (cdxi553m ^ cdxi554m ^ cdxi555m ^ cdxi556m ^ cdxi557m ^ cdxi558m ^ cdxi552m);
wire cdxi560m = reg_0_0&cdxi559m;
wire cdxi561m = cdxi504m&cdxi207m ^ r49m;
wire cdxi562m = cdxi196m&cdxi207m;
wire cdxi563m = cdxi219m&cdxi207m;
wire cdxi564m = cdxi196m&cdxi271m;
wire cdxi565m = cdxi219m&cdxi325m;
wire cdxi566m = cdxi219m&cdxi326m;
wire cdxi567m = cdxi207m&r14m;
wire cdxi568m = cdxi196m&r17m;
wire cdxi569m = cdxi219m&r24m;
wire cdxi570m = (cdxi561m ^ cdxi564m ^ cdxi565m ^ cdxi566m ^ cdxi567m ^ cdxi568m ^ cdxi569m);
wire cdxi571m = a0&cdxi570m;
wire cdxi572m = (reg_0_57);
wire cdxi573m = reg_0_4&cdxi276m;
wire cdxi574m = reg_0_2&cdxi330m;
wire cdxi575m = reg_0_2&cdxi331m;
wire cdxi576m = reg_0_7&cdxi513m;
wire cdxi577m = reg_0_4&cdxi275m;
wire cdxi578m = reg_0_2&cdxi329m;
wire cdxi579m = (cdxi573m ^ cdxi574m ^ cdxi575m ^ cdxi576m ^ cdxi577m ^ cdxi578m ^ cdxi572m);
wire cdxi580m = reg_0_0&cdxi579m;
wire cdxi581m = cdxi405m&cdxi240m ^ r53m;
wire cdxi582m = cdxi184m&cdxi240m;
wire cdxi583m = cdxi196m&cdxi311m;
wire cdxi584m = cdxi184m&cdxi241m;
wire cdxi585m = cdxi184m&cdxi242m;
wire cdxi586m = cdxi240m&r18m;
wire cdxi587m = cdxi196m&r19m;
wire cdxi588m = cdxi184m&r22m;
wire cdxi589m = (cdxi581m ^ cdxi583m ^ cdxi584m ^ cdxi585m ^ cdxi586m ^ cdxi587m ^ cdxi588m);
wire cdxi590m = a0&cdxi589m;
wire cdxi591m = (reg_0_61);
wire cdxi592m = reg_0_4&cdxi316m;
wire cdxi593m = reg_0_3&cdxi246m;
wire cdxi594m = reg_0_3&cdxi247m;
wire cdxi595m = reg_0_5&cdxi285m;
wire cdxi596m = reg_0_4&cdxi315m;
wire cdxi597m = reg_0_3&cdxi245m;
wire cdxi598m = (cdxi592m ^ cdxi593m ^ cdxi594m ^ cdxi595m ^ cdxi596m ^ cdxi597m ^ cdxi591m);
wire cdxi599m = reg_0_0&cdxi598m;
wire cdxi600m = cdxi405m&cdxi218m ^ r54m;
wire cdxi601m = cdxi184m&cdxi218m;
wire cdxi602m = cdxi196m&cdxi291m;
wire cdxi603m = cdxi184m&cdxi301m;
wire cdxi604m = cdxi184m&cdxi302m;
wire cdxi605m = cdxi218m&r18m;
wire cdxi606m = cdxi196m&r20m;
wire cdxi607m = cdxi184m&r23m;
wire cdxi608m = (cdxi600m ^ cdxi602m ^ cdxi603m ^ cdxi604m ^ cdxi605m ^ cdxi606m ^ cdxi607m);
wire cdxi609m = a0&cdxi608m;
wire cdxi610m = (reg_0_62);
wire cdxi611m = reg_0_4&cdxi296m;
wire cdxi612m = reg_0_3&cdxi306m;
wire cdxi613m = reg_0_3&cdxi307m;
wire cdxi614m = reg_0_6&cdxi285m;
wire cdxi615m = reg_0_4&cdxi295m;
wire cdxi616m = reg_0_3&cdxi305m;
wire cdxi617m = (cdxi611m ^ cdxi612m ^ cdxi613m ^ cdxi614m ^ cdxi615m ^ cdxi616m ^ cdxi610m);
wire cdxi618m = reg_0_0&cdxi617m;
wire cdxi619m = cdxi184m&cdxi485m ^ r57m;
wire cdxi620m = cdxi240m&cdxi230m;
wire cdxi621m = cdxi184m&cdxi261m;
wire cdxi622m = cdxi184m&cdxi262m;
wire cdxi623m = cdxi207m&r19m;
wire cdxi624m = cdxi240m&r21m;
wire cdxi625m = cdxi184m&r26m;
wire cdxi626m = (cdxi619m ^ cdxi620m ^ cdxi621m ^ cdxi622m ^ cdxi623m ^ cdxi624m ^ cdxi625m);
wire cdxi627m = a0&cdxi626m;
wire cdxi628m = (reg_0_65);
wire cdxi629m = reg_0_5&cdxi235m;
wire cdxi630m = reg_0_3&cdxi266m;
wire cdxi631m = reg_0_3&cdxi267m;
wire cdxi632m = reg_0_7&cdxi315m;
wire cdxi633m = reg_0_5&cdxi234m;
wire cdxi634m = reg_0_3&cdxi265m;
wire cdxi635m = (cdxi629m ^ cdxi630m ^ cdxi631m ^ cdxi632m ^ cdxi633m ^ cdxi634m ^ cdxi628m);
wire cdxi636m = reg_0_0&cdxi635m;
wire cdxi637m = cdxi445m&cdxi218m ^ r59m;
wire cdxi638m = cdxi240m&cdxi218m;
wire cdxi639m = cdxi240m&cdxi301m;
wire cdxi640m = cdxi196m&cdxi251m;
wire cdxi641m = cdxi196m&cdxi252m;
wire cdxi642m = cdxi218m&r22m;
wire cdxi643m = cdxi240m&r23m;
wire cdxi644m = cdxi196m&r25m;
wire cdxi645m = (cdxi637m ^ cdxi639m ^ cdxi640m ^ cdxi641m ^ cdxi642m ^ cdxi643m ^ cdxi644m);
wire cdxi646m = a0&cdxi645m;
wire cdxi647m = (reg_0_67);
wire cdxi648m = reg_0_5&cdxi306m;
wire cdxi649m = reg_0_4&cdxi256m;
wire cdxi650m = reg_0_4&cdxi257m;
wire cdxi651m = reg_0_6&cdxi245m;
wire cdxi652m = reg_0_5&cdxi305m;
wire cdxi653m = reg_0_4&cdxi255m;
wire cdxi654m = (cdxi648m ^ cdxi649m ^ cdxi650m ^ cdxi651m ^ cdxi652m ^ cdxi653m ^ cdxi647m);
wire cdxi655m = reg_0_0&cdxi654m;
wire cdxi656m = cdxi638m&cdxi207m ^ r62m;
wire cdxi657m = cdxi218m&cdxi207m;
wire cdxi658m = cdxi218m&cdxi261m;
wire cdxi659m = cdxi240m&cdxi337m;
wire cdxi660m = cdxi240m&cdxi338m;
wire cdxi661m = cdxi207m&r25m;
wire cdxi662m = cdxi218m&r26m;
wire cdxi663m = cdxi240m&r27m;
wire cdxi664m = (cdxi656m ^ cdxi658m ^ cdxi659m ^ cdxi660m ^ cdxi661m ^ cdxi662m ^ cdxi663m);
wire cdxi665m = a0&cdxi664m;
wire cdxi666m = (reg_0_70);
wire cdxi667m = reg_0_6&cdxi266m;
wire cdxi668m = reg_0_5&cdxi342m;
wire cdxi669m = reg_0_5&cdxi343m;
wire cdxi670m = reg_0_7&cdxi255m;
wire cdxi671m = reg_0_6&cdxi265m;
wire cdxi672m = reg_0_5&cdxi341m;
wire cdxi673m = (cdxi667m ^ cdxi668m ^ cdxi669m ^ cdxi670m ^ cdxi671m ^ cdxi672m ^ cdxi666m);
wire cdxi674m = reg_0_0&cdxi673m;
wire cdxi675m = cdxi361m&cdxi240m ^ r44m;
wire cdxi676m = cdxi582m&r1m;
wire cdxi677m = cdxi219m&cdxi311m;
wire cdxi678m = cdxi219m&cdxi312m;
wire cdxi679m = cdxi240m&r13m;
wire cdxi680m = cdxi184m&r15m;
wire cdxi681m = cdxi219m&r19m;
wire cdxi682m = (cdxi675m ^ cdxi676m ^ cdxi677m ^ cdxi678m ^ cdxi679m ^ cdxi680m ^ cdxi681m);
wire cdxi683m = cdxi185m&cdxi682m;
wire cdxi684m = (reg_0_52);
wire cdxi685m = reg_0_3&reg_0_5&cdxi136m;
wire cdxi686m = reg_0_2&cdxi316m;
wire cdxi687m = reg_0_2&cdxi317m;
wire cdxi688m = reg_0_5&cdxi373m;
wire cdxi689m = reg_0_3&cdxi533m;
wire cdxi690m = reg_0_2&cdxi315m;
wire cdxi691m = (cdxi685m ^ cdxi686m ^ cdxi687m ^ cdxi688m ^ cdxi689m ^ cdxi690m ^ cdxi684m);
wire cdxi692m = reg_0_1&cdxi691m;
wire cdxi693m = cdxi361m&cdxi218m ^ r45m;
wire cdxi694m = cdxi184m&cdxi220m;
wire cdxi695m = cdxi219m&cdxi291m;
wire cdxi696m = cdxi219m&cdxi292m;
wire cdxi697m = cdxi218m&r13m;
wire cdxi698m = cdxi184m&r16m;
wire cdxi699m = cdxi219m&r20m;
wire cdxi700m = (cdxi693m ^ cdxi694m ^ cdxi695m ^ cdxi696m ^ cdxi697m ^ cdxi698m ^ cdxi699m);
wire cdxi701m = cdxi185m&cdxi700m;
wire cdxi702m = (reg_0_53);
wire cdxi703m = reg_0_3&cdxi225m;
wire cdxi704m = reg_0_2&cdxi296m;
wire cdxi705m = reg_0_2&cdxi297m;
wire cdxi706m = reg_0_6&cdxi373m;
wire cdxi707m = reg_0_3&cdxi224m;
wire cdxi708m = reg_0_2&cdxi295m;
wire cdxi709m = (cdxi703m ^ cdxi704m ^ cdxi705m ^ cdxi706m ^ cdxi707m ^ cdxi708m ^ cdxi702m);
wire cdxi710m = reg_0_1&cdxi709m;
wire cdxi711m = cdxi185m&cdxi550m;
wire cdxi712m = reg_0_1&cdxi559m;
wire cdxi713m = cdxi185m&cdxi570m;
wire cdxi714m = reg_0_1&cdxi579m;
wire cdxi715m = cdxi524m&cdxi218m ^ r50m;
wire cdxi716m = cdxi240m&cdxi220m;
wire cdxi717m = cdxi219m&cdxi251m;
wire cdxi718m = cdxi219m&cdxi252m;
wire cdxi719m = cdxi218m&r15m;
wire cdxi720m = cdxi240m&r16m;
wire cdxi721m = cdxi219m&r25m;
wire cdxi722m = (cdxi715m ^ cdxi716m ^ cdxi717m ^ cdxi718m ^ cdxi719m ^ cdxi720m ^ cdxi721m);
wire cdxi723m = cdxi185m&cdxi722m;
wire cdxi724m = (reg_0_58);
wire cdxi725m = reg_0_5&cdxi225m;
wire cdxi726m = reg_0_2&cdxi256m;
wire cdxi727m = reg_0_2&cdxi257m;
wire cdxi728m = reg_0_6&cdxi533m;
wire cdxi729m = reg_0_5&cdxi224m;
wire cdxi730m = reg_0_2&cdxi255m;
wire cdxi731m = (cdxi725m ^ cdxi726m ^ cdxi727m ^ cdxi728m ^ cdxi729m ^ cdxi730m ^ cdxi724m);
wire cdxi732m = reg_0_1&cdxi731m;
wire cdxi733m = cdxi219m&cdxi485m ^ r51m;
wire cdxi734m = cdxi240m&cdxi271m;
wire cdxi735m = cdxi219m&cdxi261m;
wire cdxi736m = cdxi219m&cdxi262m;
wire cdxi737m = cdxi207m&r15m;
wire cdxi738m = cdxi240m&r17m;
wire cdxi739m = cdxi219m&r26m;
wire cdxi740m = (cdxi733m ^ cdxi734m ^ cdxi735m ^ cdxi736m ^ cdxi737m ^ cdxi738m ^ cdxi739m);
wire cdxi741m = cdxi185m&cdxi740m;
wire cdxi742m = (reg_0_59);
wire cdxi743m = reg_0_5&cdxi276m;
wire cdxi744m = reg_0_2&cdxi266m;
wire cdxi745m = reg_0_2&cdxi267m;
wire cdxi746m = reg_0_7&cdxi533m;
wire cdxi747m = reg_0_5&cdxi275m;
wire cdxi748m = reg_0_2&cdxi265m;
wire cdxi749m = (cdxi743m ^ cdxi744m ^ cdxi745m ^ cdxi746m ^ cdxi747m ^ cdxi748m ^ cdxi742m);
wire cdxi750m = reg_0_1&cdxi749m;
wire cdxi751m = cdxi185m&cdxi589m;
wire cdxi752m = reg_0_1&cdxi598m;
wire cdxi753m = cdxi185m&cdxi626m;
wire cdxi754m = reg_0_1&cdxi635m;
wire cdxi755m = cdxi185m&cdxi645m;
wire cdxi756m = reg_0_1&cdxi654m;
wire cdxi757m = cdxi466m&cdxi207m ^ r61m;
wire cdxi758m = cdxi218m&cdxi325m;
wire cdxi759m = cdxi196m&cdxi337m;
wire cdxi760m = cdxi196m&cdxi338m;
wire cdxi761m = cdxi207m&r23m;
wire cdxi762m = cdxi218m&r24m;
wire cdxi763m = cdxi196m&r27m;
wire cdxi764m = (cdxi757m ^ cdxi758m ^ cdxi759m ^ cdxi760m ^ cdxi761m ^ cdxi762m ^ cdxi763m);
wire cdxi765m = cdxi185m&cdxi764m;
wire cdxi766m = (reg_0_69);
wire cdxi767m = reg_0_6&cdxi330m;
wire cdxi768m = reg_0_4&cdxi342m;
wire cdxi769m = reg_0_4&cdxi343m;
wire cdxi770m = reg_0_7&cdxi305m;
wire cdxi771m = reg_0_6&cdxi329m;
wire cdxi772m = reg_0_4&cdxi341m;
wire cdxi773m = (cdxi767m ^ cdxi768m ^ cdxi769m ^ cdxi770m ^ cdxi771m ^ cdxi772m ^ cdxi766m);
wire cdxi774m = reg_0_1&cdxi773m;
wire cdxi775m = cdxi219m&cdxi589m;
wire cdxi776m = reg_0_2&cdxi598m;
wire cdxi777m = cdxi405m&cdxi207m ^ r55m;
wire cdxi778m = cdxi196m&cdxi230m;
wire cdxi779m = cdxi184m&cdxi325m;
wire cdxi780m = cdxi184m&cdxi326m;
wire cdxi781m = cdxi207m&r18m;
wire cdxi782m = cdxi196m&r21m;
wire cdxi783m = cdxi184m&r24m;
wire cdxi784m = (cdxi777m ^ cdxi778m ^ cdxi779m ^ cdxi780m ^ cdxi781m ^ cdxi782m ^ cdxi783m);
wire cdxi785m = cdxi219m&cdxi784m;
wire cdxi786m = (reg_0_63);
wire cdxi787m = reg_0_4&cdxi235m;
wire cdxi788m = reg_0_3&cdxi330m;
wire cdxi789m = reg_0_3&cdxi331m;
wire cdxi790m = reg_0_7&cdxi285m;
wire cdxi791m = reg_0_4&cdxi234m;
wire cdxi792m = reg_0_3&cdxi329m;
wire cdxi793m = (cdxi787m ^ cdxi788m ^ cdxi789m ^ cdxi790m ^ cdxi791m ^ cdxi792m ^ cdxi786m);
wire cdxi794m = reg_0_2&cdxi793m;
wire cdxi795m = cdxi219m&cdxi626m;
wire cdxi796m = reg_0_2&cdxi635m;
wire cdxi797m = cdxi219m&cdxi664m;
wire cdxi798m = reg_0_2&cdxi673m;
wire cdxi799m = cdxi184m&cdxi645m;
wire cdxi800m = reg_0_3&cdxi654m;
wire cdxi801m = cdxi445m&cdxi207m ^ r60m;
wire cdxi802m = cdxi240m&cdxi325m;
wire cdxi803m = cdxi196m&cdxi261m;
wire cdxi804m = cdxi196m&cdxi262m;
wire cdxi805m = cdxi207m&r22m;
wire cdxi806m = cdxi240m&r24m;
wire cdxi807m = cdxi196m&r26m;
wire cdxi808m = (cdxi801m ^ cdxi802m ^ cdxi803m ^ cdxi804m ^ cdxi805m ^ cdxi806m ^ cdxi807m);
wire cdxi809m = cdxi184m&cdxi808m;
wire cdxi810m = (reg_0_68);
wire cdxi811m = reg_0_5&cdxi330m;
wire cdxi812m = reg_0_4&cdxi266m;
wire cdxi813m = reg_0_4&cdxi267m;
wire cdxi814m = reg_0_7&cdxi245m;
wire cdxi815m = reg_0_5&cdxi329m;
wire cdxi816m = reg_0_4&cdxi265m;
wire cdxi817m = (cdxi811m ^ cdxi812m ^ cdxi813m ^ cdxi814m ^ cdxi815m ^ cdxi816m ^ cdxi810m);
wire cdxi818m = reg_0_3&cdxi817m;
wire cdxi819m = cdxi184m&cdxi764m;
wire cdxi820m = reg_0_3&cdxi773m;
wire cdxi821m = cdxi185m&cdxi361m&cdxi196m ^ r63m;
wire cdxi822m = cdxi361m&cdxi196m;
wire cdxi823m = cdxi362m&cdxi196m;
wire cdxi824m = cdxi363m&cdxi196m;
wire cdxi825m = cdxi185m&cdxi361m;
wire cdxi826m = cdxi361m&cdxi197m;
wire cdxi827m = cdxi823m&r1m;
wire cdxi828m = cdxi363m&cdxi281m;
wire cdxi829m = cdxi363m&cdxi282m;
wire cdxi830m = cdxi405m&r7m;
wire cdxi831m = cdxi219m&cdxi410m;
wire cdxi832m = cdxi361m&r9m;
wire cdxi833m = cdxi406m&r13m;
wire cdxi834m = cdxi362m&r14m;
wire cdxi835m = cdxi363m&r18m;
wire cdxi836m = cdxi196m&r28m;
wire cdxi837m = cdxi184m&r29m;
wire cdxi838m = cdxi219m&r33m;
wire cdxi839m = cdxi185m&r43m;
wire cdxi840m = (cdxi821m ^ cdxi826m ^ cdxi827m ^ cdxi828m ^ cdxi829m ^ cdxi830m ^ cdxi831m ^ cdxi832m ^ cdxi833m ^ cdxi834m ^ cdxi835m ^ cdxi836m ^ cdxi837m ^ cdxi838m ^ cdxi839m);
wire cdxi841m = a0&cdxi840m;
wire cdxi842m = (reg_0_37);
wire cdxi843m = (reg_0_71);
wire cdxi844m = reg_0_2&cdxi416m;
wire cdxi845m = reg_0_1&cdxi515m;
wire cdxi846m = reg_0_1&cdxi516m;
wire cdxi847m = reg_0_1&cdxi517m;
wire cdxi848m = reg_0_3&reg_0_4&cdxi372m;
wire cdxi849m = reg_0_2&cdxi419m;
wire cdxi850m = reg_0_2&cdxi420m;
wire cdxi851m = reg_0_1&cdxi518m;
wire cdxi852m = reg_0_1&cdxi519m;
wire cdxi853m = reg_0_1&cdxi520m;
wire cdxi854m = reg_0_4&cdxi374m;
wire cdxi855m = reg_0_3&cdxi842m;
wire cdxi856m = reg_0_2&cdxi415m;
wire cdxi857m = reg_0_1&cdxi514m;
wire cdxi858m = (cdxi844m ^ cdxi845m ^ cdxi846m ^ cdxi847m ^ cdxi848m ^ cdxi849m ^ cdxi850m ^ cdxi851m ^ cdxi852m ^ cdxi853m ^ cdxi854m ^ cdxi855m ^ cdxi856m ^ cdxi857m ^ cdxi843m);
wire cdxi859m = reg_0_0&cdxi858m;
wire cdxi860m = cdxi825m&cdxi240m ^ r64m;
wire cdxi861m = cdxi361m&cdxi240m;
wire cdxi862m = cdxi362m&cdxi240m;
wire cdxi863m = cdxi363m&cdxi240m;
wire cdxi864m = cdxi861m&r0m;
wire cdxi865m = cdxi862m&r1m;
wire cdxi866m = cdxi363m&cdxi311m;
wire cdxi867m = cdxi363m&cdxi312m;
wire cdxi868m = cdxi582m&r7m;
wire cdxi869m = cdxi524m&r8m;
wire cdxi870m = cdxi361m&r10m;
wire cdxi871m = cdxi446m&r13m;
wire cdxi872m = cdxi362m&r15m;
wire cdxi873m = cdxi363m&r19m;
wire cdxi874m = cdxi240m&r28m;
wire cdxi875m = cdxi184m&r30m;
wire cdxi876m = cdxi219m&r34m;
wire cdxi877m = cdxi185m&r44m;
wire cdxi878m = (cdxi860m ^ cdxi864m ^ cdxi865m ^ cdxi866m ^ cdxi867m ^ cdxi868m ^ cdxi869m ^ cdxi870m ^ cdxi871m ^ cdxi872m ^ cdxi873m ^ cdxi874m ^ cdxi875m ^ cdxi876m ^ cdxi877m);
wire cdxi879m = a0&cdxi878m;
wire cdxi880m = (reg_0_38);
wire cdxi881m = (reg_0_42);
wire cdxi882m = (reg_0_72);
wire cdxi883m = reg_0_2&reg_0_3&reg_0_5&cdxi130m;
wire cdxi884m = reg_0_1&cdxi685m;
wire cdxi885m = reg_0_1&cdxi686m;
wire cdxi886m = reg_0_1&cdxi687m;
wire cdxi887m = reg_0_3&reg_0_5&cdxi372m;
wire cdxi888m = reg_0_2&reg_0_5&cdxi190m;
wire cdxi889m = reg_0_2&reg_0_3&cdxi455m;
wire cdxi890m = reg_0_1&cdxi688m;
wire cdxi891m = reg_0_1&cdxi689m;
wire cdxi892m = reg_0_1&cdxi690m;
wire cdxi893m = reg_0_5&cdxi374m;
wire cdxi894m = reg_0_3&cdxi880m;
wire cdxi895m = reg_0_2&cdxi881m;
wire cdxi896m = reg_0_1&cdxi684m;
wire cdxi897m = (cdxi883m ^ cdxi884m ^ cdxi885m ^ cdxi886m ^ cdxi887m ^ cdxi888m ^ cdxi889m ^ cdxi890m ^ cdxi891m ^ cdxi892m ^ cdxi893m ^ cdxi894m ^ cdxi895m ^ cdxi896m ^ cdxi882m);
wire cdxi898m = reg_0_0&cdxi897m;
wire cdxi899m = cdxi825m&cdxi218m ^ r65m;
wire cdxi900m = cdxi361m&cdxi218m;
wire cdxi901m = cdxi362m&cdxi218m;
wire cdxi902m = cdxi363m&cdxi218m;
wire cdxi903m = cdxi900m&r0m;
wire cdxi904m = cdxi362m&cdxi220m;
wire cdxi905m = cdxi363m&cdxi291m;
wire cdxi906m = cdxi363m&cdxi292m;
wire cdxi907m = cdxi184m&cdxi389m;
wire cdxi908m = cdxi384m&r8m;
wire cdxi909m = cdxi361m&r11m;
wire cdxi910m = cdxi385m&r13m;
wire cdxi911m = cdxi362m&r16m;
wire cdxi912m = cdxi363m&r20m;
wire cdxi913m = cdxi218m&r28m;
wire cdxi914m = cdxi184m&r31m;
wire cdxi915m = cdxi219m&r35m;
wire cdxi916m = cdxi185m&r45m;
wire cdxi917m = (cdxi899m ^ cdxi903m ^ cdxi904m ^ cdxi905m ^ cdxi906m ^ cdxi907m ^ cdxi908m ^ cdxi909m ^ cdxi910m ^ cdxi911m ^ cdxi912m ^ cdxi913m ^ cdxi914m ^ cdxi915m ^ cdxi916m);
wire cdxi918m = a0&cdxi917m;
wire cdxi919m = (reg_0_43);
wire cdxi920m = (reg_0_73);
wire cdxi921m = reg_0_2&reg_0_3&reg_0_6&cdxi130m;
wire cdxi922m = reg_0_1&cdxi703m;
wire cdxi923m = reg_0_1&cdxi704m;
wire cdxi924m = reg_0_1&cdxi705m;
wire cdxi925m = reg_0_3&cdxi399m;
wire cdxi926m = reg_0_2&reg_0_6&cdxi190m;
wire cdxi927m = reg_0_2&reg_0_3&cdxi394m;
wire cdxi928m = reg_0_1&cdxi706m;
wire cdxi929m = reg_0_1&cdxi707m;
wire cdxi930m = reg_0_1&cdxi708m;
wire cdxi931m = reg_0_6&cdxi374m;
wire cdxi932m = reg_0_3&cdxi395m;
wire cdxi933m = reg_0_2&cdxi919m;
wire cdxi934m = reg_0_1&cdxi702m;
wire cdxi935m = (cdxi921m ^ cdxi922m ^ cdxi923m ^ cdxi924m ^ cdxi925m ^ cdxi926m ^ cdxi927m ^ cdxi928m ^ cdxi929m ^ cdxi930m ^ cdxi931m ^ cdxi932m ^ cdxi933m ^ cdxi934m ^ cdxi920m);
wire cdxi936m = reg_0_0&cdxi935m;
wire cdxi937m = cdxi825m&cdxi207m ^ r66m;
wire cdxi938m = cdxi361m&cdxi207m;
wire cdxi939m = cdxi362m&cdxi207m;
wire cdxi940m = cdxi363m&cdxi207m;
wire cdxi941m = cdxi361m&cdxi208m;
wire cdxi942m = cdxi362m&cdxi271m;
wire cdxi943m = cdxi363m&cdxi230m;
wire cdxi944m = cdxi363m&cdxi231m;
wire cdxi945m = cdxi425m&r7m;
wire cdxi946m = cdxi219m&cdxi430m;
wire cdxi947m = cdxi361m&r12m;
wire cdxi948m = cdxi426m&r13m;
wire cdxi949m = cdxi362m&r17m;
wire cdxi950m = cdxi363m&r21m;
wire cdxi951m = cdxi207m&r28m;
wire cdxi952m = cdxi184m&r32m;
wire cdxi953m = cdxi219m&r36m;
wire cdxi954m = cdxi185m&r46m;
wire cdxi955m = (cdxi937m ^ cdxi941m ^ cdxi942m ^ cdxi943m ^ cdxi944m ^ cdxi945m ^ cdxi946m ^ cdxi947m ^ cdxi948m ^ cdxi949m ^ cdxi950m ^ cdxi951m ^ cdxi952m ^ cdxi953m ^ cdxi954m);
wire cdxi956m = a0&cdxi955m;
wire cdxi957m = (reg_0_40);
wire cdxi958m = (reg_0_54);
wire cdxi959m = (reg_0_74);
wire cdxi960m = reg_0_2&cdxi436m;
wire cdxi961m = reg_0_1&reg_0_3&cdxi276m;
wire cdxi962m = reg_0_1&reg_0_2&cdxi235m;
wire cdxi963m = reg_0_1&reg_0_2&cdxi236m;
wire cdxi964m = reg_0_3&reg_0_7&cdxi372m;
wire cdxi965m = reg_0_2&cdxi439m;
wire cdxi966m = reg_0_2&cdxi440m;
wire cdxi967m = reg_0_1&reg_0_7&cdxi373m;
wire cdxi968m = reg_0_1&reg_0_3&cdxi275m;
wire cdxi969m = reg_0_1&reg_0_2&cdxi234m;
wire cdxi970m = reg_0_7&cdxi374m;
wire cdxi971m = reg_0_3&cdxi957m;
wire cdxi972m = reg_0_2&cdxi435m;
wire cdxi973m = reg_0_1&cdxi958m;
wire cdxi974m = (cdxi960m ^ cdxi961m ^ cdxi962m ^ cdxi963m ^ cdxi964m ^ cdxi965m ^ cdxi966m ^ cdxi967m ^ cdxi968m ^ cdxi969m ^ cdxi970m ^ cdxi971m ^ cdxi972m ^ cdxi973m ^ cdxi959m);
wire cdxi975m = reg_0_0&cdxi974m;
wire cdxi976m = cdxi363m&cdxi466m ^ r68m;
wire cdxi977m = cdxi219m&cdxi466m;
wire cdxi978m = cdxi406m&cdxi218m;
wire cdxi979m = cdxi219m&cdxi467m;
wire cdxi980m = cdxi406m&cdxi220m;
wire cdxi981m = cdxi363m&cdxi301m;
wire cdxi982m = cdxi363m&cdxi302m;
wire cdxi983m = cdxi196m&cdxi389m;
wire cdxi984m = cdxi384m&r9m;
wire cdxi985m = cdxi219m&cdxi471m;
wire cdxi986m = cdxi385m&r14m;
wire cdxi987m = cdxi406m&r16m;
wire cdxi988m = cdxi363m&r23m;
wire cdxi989m = cdxi218m&r29m;
wire cdxi990m = cdxi196m&r31m;
wire cdxi991m = cdxi219m&r38m;
wire cdxi992m = cdxi185m&r48m;
wire cdxi993m = (cdxi976m ^ cdxi979m ^ cdxi980m ^ cdxi981m ^ cdxi982m ^ cdxi983m ^ cdxi984m ^ cdxi985m ^ cdxi986m ^ cdxi987m ^ cdxi988m ^ cdxi989m ^ cdxi990m ^ cdxi991m ^ cdxi992m);
wire cdxi994m = a0&cdxi993m;
wire cdxi995m = (reg_0_76);
wire cdxi996m = reg_0_2&cdxi476m;
wire cdxi997m = reg_0_1&cdxi553m;
wire cdxi998m = reg_0_1&cdxi554m;
wire cdxi999m = reg_0_1&cdxi555m;
wire cdxi1000m = reg_0_4&cdxi399m;
wire cdxi1001m = reg_0_2&cdxi479m;
wire cdxi1002m = reg_0_2&cdxi480m;
wire cdxi1003m = reg_0_1&cdxi556m;
wire cdxi1004m = reg_0_1&cdxi557m;
wire cdxi1005m = reg_0_1&cdxi558m;
wire cdxi1006m = reg_0_6&cdxi842m;
wire cdxi1007m = reg_0_4&cdxi395m;
wire cdxi1008m = reg_0_2&cdxi475m;
wire cdxi1009m = reg_0_1&cdxi552m;
wire cdxi1010m = (cdxi996m ^ cdxi997m ^ cdxi998m ^ cdxi999m ^ cdxi1000m ^ cdxi1001m ^ cdxi1002m ^ cdxi1003m ^ cdxi1004m ^ cdxi1005m ^ cdxi1006m ^ cdxi1007m ^ cdxi1008m ^ cdxi1009m ^ cdxi995m);
wire cdxi1011m = reg_0_0&cdxi1010m;
wire cdxi1012m = cdxi363m&cdxi638m ^ r70m;
wire cdxi1013m = cdxi524m&cdxi218m;
wire cdxi1014m = cdxi446m&cdxi218m;
wire cdxi1015m = cdxi1013m&r0m;
wire cdxi1016m = cdxi446m&cdxi220m;
wire cdxi1017m = cdxi363m&cdxi251m;
wire cdxi1018m = cdxi363m&cdxi252m;
wire cdxi1019m = cdxi240m&cdxi389m;
wire cdxi1020m = cdxi384m&r10m;
wire cdxi1021m = cdxi524m&r11m;
wire cdxi1022m = cdxi385m&r15m;
wire cdxi1023m = cdxi446m&r16m;
wire cdxi1024m = cdxi363m&r25m;
wire cdxi1025m = cdxi218m&r30m;
wire cdxi1026m = cdxi240m&r31m;
wire cdxi1027m = cdxi219m&r40m;
wire cdxi1028m = cdxi185m&r50m;
wire cdxi1029m = (cdxi1012m ^ cdxi1015m ^ cdxi1016m ^ cdxi1017m ^ cdxi1018m ^ cdxi1019m ^ cdxi1020m ^ cdxi1021m ^ cdxi1022m ^ cdxi1023m ^ cdxi1024m ^ cdxi1025m ^ cdxi1026m ^ cdxi1027m ^ cdxi1028m);
wire cdxi1030m = a0&cdxi1029m;
wire cdxi1031m = (reg_0_48);
wire cdxi1032m = (reg_0_78);
wire cdxi1033m = reg_0_2&reg_0_5&reg_0_6&cdxi130m;
wire cdxi1034m = reg_0_1&cdxi725m;
wire cdxi1035m = reg_0_1&cdxi726m;
wire cdxi1036m = reg_0_1&cdxi727m;
wire cdxi1037m = reg_0_5&cdxi399m;
wire cdxi1038m = reg_0_2&reg_0_6&cdxi455m;
wire cdxi1039m = reg_0_2&reg_0_5&cdxi394m;
wire cdxi1040m = reg_0_1&cdxi728m;
wire cdxi1041m = reg_0_1&cdxi729m;
wire cdxi1042m = reg_0_1&cdxi730m;
wire cdxi1043m = reg_0_6&cdxi880m;
wire cdxi1044m = reg_0_5&cdxi395m;
wire cdxi1045m = reg_0_2&cdxi1031m;
wire cdxi1046m = reg_0_1&cdxi724m;
wire cdxi1047m = (cdxi1033m ^ cdxi1034m ^ cdxi1035m ^ cdxi1036m ^ cdxi1037m ^ cdxi1038m ^ cdxi1039m ^ cdxi1040m ^ cdxi1041m ^ cdxi1042m ^ cdxi1043m ^ cdxi1044m ^ cdxi1045m ^ cdxi1046m ^ cdxi1032m);
wire cdxi1048m = reg_0_0&cdxi1047m;
wire cdxi1049m = cdxi363m&cdxi657m ^ r72m;
wire cdxi1050m = cdxi384m&cdxi207m;
wire cdxi1051m = cdxi385m&cdxi207m;
wire cdxi1052m = cdxi384m&cdxi208m;
wire cdxi1053m = cdxi385m&cdxi271m;
wire cdxi1054m = cdxi363m&cdxi337m;
wire cdxi1055m = cdxi363m&cdxi338m;
wire cdxi1056m = cdxi657m&r7m;
wire cdxi1057m = cdxi563m&r11m;
wire cdxi1058m = cdxi384m&r12m;
wire cdxi1059m = cdxi426m&r16m;
wire cdxi1060m = cdxi385m&r17m;
wire cdxi1061m = cdxi363m&r27m;
wire cdxi1062m = cdxi207m&r31m;
wire cdxi1063m = cdxi218m&r32m;
wire cdxi1064m = cdxi219m&r42m;
wire cdxi1065m = cdxi185m&r52m;
wire cdxi1066m = (cdxi1049m ^ cdxi1052m ^ cdxi1053m ^ cdxi1054m ^ cdxi1055m ^ cdxi1056m ^ cdxi1057m ^ cdxi1058m ^ cdxi1059m ^ cdxi1060m ^ cdxi1061m ^ cdxi1062m ^ cdxi1063m ^ cdxi1064m ^ cdxi1065m);
wire cdxi1067m = a0&cdxi1066m;
wire cdxi1068m = (reg_0_50);
wire cdxi1069m = (reg_0_60);
wire cdxi1070m = (reg_0_80);
wire cdxi1071m = reg_0_2&reg_0_6&cdxi213m;
wire cdxi1072m = reg_0_1&reg_0_6&cdxi276m;
wire cdxi1073m = reg_0_1&reg_0_2&cdxi342m;
wire cdxi1074m = reg_0_1&reg_0_2&cdxi343m;
wire cdxi1075m = reg_0_6&reg_0_7&cdxi372m;
wire cdxi1076m = reg_0_2&reg_0_7&cdxi394m;
wire cdxi1077m = reg_0_2&reg_0_6&cdxi212m;
wire cdxi1078m = reg_0_1&reg_0_7&cdxi224m;
wire cdxi1079m = reg_0_1&reg_0_6&cdxi275m;
wire cdxi1080m = reg_0_1&reg_0_2&cdxi341m;
wire cdxi1081m = reg_0_7&cdxi395m;
wire cdxi1082m = reg_0_6&cdxi957m;
wire cdxi1083m = reg_0_2&cdxi1068m;
wire cdxi1084m = reg_0_1&cdxi1069m;
wire cdxi1085m = (cdxi1071m ^ cdxi1072m ^ cdxi1073m ^ cdxi1074m ^ cdxi1075m ^ cdxi1076m ^ cdxi1077m ^ cdxi1078m ^ cdxi1079m ^ cdxi1080m ^ cdxi1081m ^ cdxi1082m ^ cdxi1083m ^ cdxi1084m ^ cdxi1070m);
wire cdxi1086m = reg_0_0&cdxi1085m;
wire cdxi1087m = cdxi362m&cdxi466m ^ r74m;
wire cdxi1088m = cdxi405m&cdxi218m;
wire cdxi1089m = cdxi1088m&r0m;
wire cdxi1090m = cdxi406m&cdxi291m;
wire cdxi1091m = cdxi362m&cdxi301m;
wire cdxi1092m = cdxi362m&cdxi302m;
wire cdxi1093m = cdxi466m&r8m;
wire cdxi1094m = cdxi184m&cdxi470m;
wire cdxi1095m = cdxi405m&r11m;
wire cdxi1096m = cdxi385m&r18m;
wire cdxi1097m = cdxi406m&r20m;
wire cdxi1098m = cdxi362m&r23m;
wire cdxi1099m = cdxi218m&r33m;
wire cdxi1100m = cdxi196m&r35m;
wire cdxi1101m = cdxi184m&r38m;
wire cdxi1102m = cdxi185m&r54m;
wire cdxi1103m = (cdxi1087m ^ cdxi1089m ^ cdxi1090m ^ cdxi1091m ^ cdxi1092m ^ cdxi1093m ^ cdxi1094m ^ cdxi1095m ^ cdxi1096m ^ cdxi1097m ^ cdxi1098m ^ cdxi1099m ^ cdxi1100m ^ cdxi1101m ^ cdxi1102m);
wire cdxi1104m = a0&cdxi1103m;
wire cdxi1105m = (reg_0_82);
wire cdxi1106m = reg_0_3&cdxi476m;
wire cdxi1107m = reg_0_1&cdxi611m;
wire cdxi1108m = reg_0_1&cdxi612m;
wire cdxi1109m = reg_0_1&cdxi613m;
wire cdxi1110m = reg_0_4&reg_0_6&cdxi190m;
wire cdxi1111m = reg_0_3&cdxi479m;
wire cdxi1112m = reg_0_3&cdxi480m;
wire cdxi1113m = reg_0_1&cdxi614m;
wire cdxi1114m = reg_0_1&cdxi615m;
wire cdxi1115m = reg_0_1&cdxi616m;
wire cdxi1116m = reg_0_6&cdxi415m;
wire cdxi1117m = reg_0_4&cdxi919m;
wire cdxi1118m = reg_0_3&cdxi475m;
wire cdxi1119m = reg_0_1&cdxi610m;
wire cdxi1120m = (cdxi1106m ^ cdxi1107m ^ cdxi1108m ^ cdxi1109m ^ cdxi1110m ^ cdxi1111m ^ cdxi1112m ^ cdxi1113m ^ cdxi1114m ^ cdxi1115m ^ cdxi1116m ^ cdxi1117m ^ cdxi1118m ^ cdxi1119m ^ cdxi1105m);
wire cdxi1121m = reg_0_0&cdxi1120m;
wire cdxi1122m = cdxi362m&cdxi562m ^ r75m;
wire cdxi1123m = cdxi405m&cdxi207m;
wire cdxi1124m = cdxi406m&cdxi207m;
wire cdxi1125m = cdxi405m&cdxi208m;
wire cdxi1126m = cdxi406m&cdxi230m;
wire cdxi1127m = cdxi362m&cdxi325m;
wire cdxi1128m = cdxi362m&cdxi326m;
wire cdxi1129m = cdxi196m&cdxi430m;
wire cdxi1130m = cdxi425m&r9m;
wire cdxi1131m = cdxi405m&r12m;
wire cdxi1132m = cdxi426m&r18m;
wire cdxi1133m = cdxi406m&r21m;
wire cdxi1134m = cdxi362m&r24m;
wire cdxi1135m = cdxi207m&r33m;
wire cdxi1136m = cdxi196m&r36m;
wire cdxi1137m = cdxi184m&r39m;
wire cdxi1138m = cdxi185m&r55m;
wire cdxi1139m = (cdxi1122m ^ cdxi1125m ^ cdxi1126m ^ cdxi1127m ^ cdxi1128m ^ cdxi1129m ^ cdxi1130m ^ cdxi1131m ^ cdxi1132m ^ cdxi1133m ^ cdxi1134m ^ cdxi1135m ^ cdxi1136m ^ cdxi1137m ^ cdxi1138m);
wire cdxi1140m = a0&cdxi1139m;
wire cdxi1141m = (reg_0_47);
wire cdxi1142m = (reg_0_83);
wire cdxi1143m = reg_0_3&reg_0_4&cdxi213m;
wire cdxi1144m = reg_0_1&cdxi787m;
wire cdxi1145m = reg_0_1&cdxi788m;
wire cdxi1146m = reg_0_1&cdxi789m;
wire cdxi1147m = reg_0_4&cdxi439m;
wire cdxi1148m = reg_0_3&reg_0_7&cdxi201m;
wire cdxi1149m = reg_0_3&reg_0_4&cdxi212m;
wire cdxi1150m = reg_0_1&cdxi790m;
wire cdxi1151m = reg_0_1&cdxi791m;
wire cdxi1152m = reg_0_1&cdxi792m;
wire cdxi1153m = reg_0_7&cdxi415m;
wire cdxi1154m = reg_0_4&cdxi435m;
wire cdxi1155m = reg_0_3&cdxi1141m;
wire cdxi1156m = reg_0_1&cdxi786m;
wire cdxi1157m = (cdxi1143m ^ cdxi1144m ^ cdxi1145m ^ cdxi1146m ^ cdxi1147m ^ cdxi1148m ^ cdxi1149m ^ cdxi1150m ^ cdxi1151m ^ cdxi1152m ^ cdxi1153m ^ cdxi1154m ^ cdxi1155m ^ cdxi1156m ^ cdxi1142m);
wire cdxi1158m = reg_0_0&cdxi1157m;
wire cdxi1159m = cdxi362m&cdxi485m ^ r77m;
wire cdxi1160m = cdxi184m&cdxi485m;
wire cdxi1161m = cdxi446m&cdxi207m;
wire cdxi1162m = cdxi184m&cdxi486m;
wire cdxi1163m = cdxi446m&cdxi230m;
wire cdxi1164m = cdxi362m&cdxi261m;
wire cdxi1165m = cdxi362m&cdxi262m;
wire cdxi1166m = cdxi240m&cdxi430m;
wire cdxi1167m = cdxi425m&r10m;
wire cdxi1168m = cdxi184m&cdxi490m;
wire cdxi1169m = cdxi426m&r19m;
wire cdxi1170m = cdxi446m&r21m;
wire cdxi1171m = cdxi362m&r26m;
wire cdxi1172m = cdxi207m&r34m;
wire cdxi1173m = cdxi240m&r36m;
wire cdxi1174m = cdxi184m&r41m;
wire cdxi1175m = cdxi185m&r57m;
wire cdxi1176m = (cdxi1159m ^ cdxi1162m ^ cdxi1163m ^ cdxi1164m ^ cdxi1165m ^ cdxi1166m ^ cdxi1167m ^ cdxi1168m ^ cdxi1169m ^ cdxi1170m ^ cdxi1171m ^ cdxi1172m ^ cdxi1173m ^ cdxi1174m ^ cdxi1175m);
wire cdxi1177m = a0&cdxi1176m;
wire cdxi1178m = (reg_0_85);
wire cdxi1179m = reg_0_3&cdxi495m;
wire cdxi1180m = reg_0_1&cdxi629m;
wire cdxi1181m = reg_0_1&cdxi630m;
wire cdxi1182m = reg_0_1&cdxi631m;
wire cdxi1183m = reg_0_5&cdxi439m;
wire cdxi1184m = reg_0_3&cdxi498m;
wire cdxi1185m = reg_0_3&cdxi499m;
wire cdxi1186m = reg_0_1&cdxi632m;
wire cdxi1187m = reg_0_1&cdxi633m;
wire cdxi1188m = reg_0_1&cdxi634m;
wire cdxi1189m = reg_0_7&cdxi881m;
wire cdxi1190m = reg_0_5&cdxi435m;
wire cdxi1191m = reg_0_3&cdxi494m;
wire cdxi1192m = reg_0_1&cdxi628m;
wire cdxi1193m = (cdxi1179m ^ cdxi1180m ^ cdxi1181m ^ cdxi1182m ^ cdxi1183m ^ cdxi1184m ^ cdxi1185m ^ cdxi1186m ^ cdxi1187m ^ cdxi1188m ^ cdxi1189m ^ cdxi1190m ^ cdxi1191m ^ cdxi1192m ^ cdxi1178m);
wire cdxi1194m = reg_0_0&cdxi1193m;
wire cdxi1195m = cdxi362m&cdxi657m ^ r78m;
wire cdxi1196m = cdxi601m&cdxi207m;
wire cdxi1197m = cdxi601m&cdxi208m;
wire cdxi1198m = cdxi385m&cdxi230m;
wire cdxi1199m = cdxi362m&cdxi337m;
wire cdxi1200m = cdxi362m&cdxi338m;
wire cdxi1201m = cdxi218m&cdxi430m;
wire cdxi1202m = cdxi425m&r11m;
wire cdxi1203m = cdxi601m&r12m;
wire cdxi1204m = cdxi426m&r20m;
wire cdxi1205m = cdxi385m&r21m;
wire cdxi1206m = cdxi362m&r27m;
wire cdxi1207m = cdxi207m&r35m;
wire cdxi1208m = cdxi218m&r36m;
wire cdxi1209m = cdxi184m&r42m;
wire cdxi1210m = cdxi185m&r58m;
wire cdxi1211m = (cdxi1195m ^ cdxi1197m ^ cdxi1198m ^ cdxi1199m ^ cdxi1200m ^ cdxi1201m ^ cdxi1202m ^ cdxi1203m ^ cdxi1204m ^ cdxi1205m ^ cdxi1206m ^ cdxi1207m ^ cdxi1208m ^ cdxi1209m ^ cdxi1210m);
wire cdxi1212m = a0&cdxi1211m;
wire cdxi1213m = (reg_0_66);
wire cdxi1214m = (reg_0_86);
wire cdxi1215m = reg_0_3&reg_0_6&cdxi213m;
wire cdxi1216m = reg_0_1&reg_0_6&cdxi235m;
wire cdxi1217m = reg_0_1&reg_0_3&cdxi342m;
wire cdxi1218m = reg_0_1&reg_0_3&cdxi343m;
wire cdxi1219m = reg_0_6&cdxi439m;
wire cdxi1220m = reg_0_3&reg_0_7&cdxi394m;
wire cdxi1221m = reg_0_3&reg_0_6&cdxi212m;
wire cdxi1222m = reg_0_1&reg_0_7&cdxi295m;
wire cdxi1223m = reg_0_1&reg_0_6&cdxi234m;
wire cdxi1224m = reg_0_1&reg_0_3&cdxi341m;
wire cdxi1225m = reg_0_7&cdxi919m;
wire cdxi1226m = reg_0_6&cdxi435m;
wire cdxi1227m = reg_0_3&cdxi1068m;
wire cdxi1228m = reg_0_1&cdxi1213m;
wire cdxi1229m = (cdxi1215m ^ cdxi1216m ^ cdxi1217m ^ cdxi1218m ^ cdxi1219m ^ cdxi1220m ^ cdxi1221m ^ cdxi1222m ^ cdxi1223m ^ cdxi1224m ^ cdxi1225m ^ cdxi1226m ^ cdxi1227m ^ cdxi1228m ^ cdxi1214m);
wire cdxi1230m = reg_0_0&cdxi1229m;
wire cdxi1231m = cdxi406m&cdxi485m ^ r80m;
wire cdxi1232m = cdxi445m&cdxi207m;
wire cdxi1233m = cdxi406m&cdxi240m;
wire cdxi1234m = cdxi445m&cdxi208m;
wire cdxi1235m = cdxi446m&cdxi325m;
wire cdxi1236m = cdxi406m&cdxi261m;
wire cdxi1237m = cdxi406m&cdxi262m;
wire cdxi1238m = cdxi485m&r9m;
wire cdxi1239m = cdxi196m&cdxi489m;
wire cdxi1240m = cdxi445m&r12m;
wire cdxi1241m = cdxi426m&r22m;
wire cdxi1242m = cdxi446m&r24m;
wire cdxi1243m = cdxi406m&r26m;
wire cdxi1244m = cdxi207m&r37m;
wire cdxi1245m = cdxi240m&r39m;
wire cdxi1246m = cdxi196m&r41m;
wire cdxi1247m = cdxi185m&r60m;
wire cdxi1248m = (cdxi1231m ^ cdxi1234m ^ cdxi1235m ^ cdxi1236m ^ cdxi1237m ^ cdxi1238m ^ cdxi1239m ^ cdxi1240m ^ cdxi1241m ^ cdxi1242m ^ cdxi1243m ^ cdxi1244m ^ cdxi1245m ^ cdxi1246m ^ cdxi1247m);
wire cdxi1249m = a0&cdxi1248m;
wire cdxi1250m = (reg_0_88);
wire cdxi1251m = reg_0_4&cdxi495m;
wire cdxi1252m = reg_0_1&cdxi811m;
wire cdxi1253m = reg_0_1&cdxi812m;
wire cdxi1254m = reg_0_1&cdxi813m;
wire cdxi1255m = reg_0_5&reg_0_7&cdxi201m;
wire cdxi1256m = reg_0_4&cdxi498m;
wire cdxi1257m = reg_0_4&cdxi499m;
wire cdxi1258m = reg_0_1&cdxi814m;
wire cdxi1259m = reg_0_1&cdxi815m;
wire cdxi1260m = reg_0_1&cdxi816m;
wire cdxi1261m = reg_0_7&cdxi456m;
wire cdxi1262m = reg_0_5&cdxi1141m;
wire cdxi1263m = reg_0_4&cdxi494m;
wire cdxi1264m = reg_0_1&cdxi810m;
wire cdxi1265m = (cdxi1251m ^ cdxi1252m ^ cdxi1253m ^ cdxi1254m ^ cdxi1255m ^ cdxi1256m ^ cdxi1257m ^ cdxi1258m ^ cdxi1259m ^ cdxi1260m ^ cdxi1261m ^ cdxi1262m ^ cdxi1263m ^ cdxi1264m ^ cdxi1250m);
wire cdxi1266m = reg_0_0&cdxi1265m;
wire cdxi1267m = cdxi406m&cdxi657m ^ r81m;
wire cdxi1268m = cdxi466m&cdxi207m;
wire cdxi1269m = cdxi466m&cdxi208m;
wire cdxi1270m = cdxi385m&cdxi325m;
wire cdxi1271m = cdxi406m&cdxi337m;
wire cdxi1272m = cdxi406m&cdxi338m;
wire cdxi1273m = cdxi657m&r9m;
wire cdxi1274m = cdxi562m&r11m;
wire cdxi1275m = cdxi466m&r12m;
wire cdxi1276m = cdxi426m&r23m;
wire cdxi1277m = cdxi385m&r24m;
wire cdxi1278m = cdxi406m&r27m;
wire cdxi1279m = cdxi207m&r38m;
wire cdxi1280m = cdxi218m&r39m;
wire cdxi1281m = cdxi196m&r42m;
wire cdxi1282m = cdxi185m&r61m;
wire cdxi1283m = (cdxi1267m ^ cdxi1269m ^ cdxi1270m ^ cdxi1271m ^ cdxi1272m ^ cdxi1273m ^ cdxi1274m ^ cdxi1275m ^ cdxi1276m ^ cdxi1277m ^ cdxi1278m ^ cdxi1279m ^ cdxi1280m ^ cdxi1281m ^ cdxi1282m);
wire cdxi1284m = a0&cdxi1283m;
wire cdxi1285m = (reg_0_89);
wire cdxi1286m = reg_0_4&reg_0_6&cdxi213m;
wire cdxi1287m = reg_0_1&cdxi767m;
wire cdxi1288m = reg_0_1&cdxi768m;
wire cdxi1289m = reg_0_1&cdxi769m;
wire cdxi1290m = reg_0_6&reg_0_7&cdxi201m;
wire cdxi1291m = reg_0_4&reg_0_7&cdxi394m;
wire cdxi1292m = reg_0_4&reg_0_6&cdxi212m;
wire cdxi1293m = reg_0_1&cdxi770m;
wire cdxi1294m = reg_0_1&cdxi771m;
wire cdxi1295m = reg_0_1&cdxi772m;
wire cdxi1296m = reg_0_7&cdxi475m;
wire cdxi1297m = reg_0_6&cdxi1141m;
wire cdxi1298m = reg_0_4&cdxi1068m;
wire cdxi1299m = reg_0_1&cdxi766m;
wire cdxi1300m = (cdxi1286m ^ cdxi1287m ^ cdxi1288m ^ cdxi1289m ^ cdxi1290m ^ cdxi1291m ^ cdxi1292m ^ cdxi1293m ^ cdxi1294m ^ cdxi1295m ^ cdxi1296m ^ cdxi1297m ^ cdxi1298m ^ cdxi1299m ^ cdxi1285m);
wire cdxi1301m = reg_0_0&cdxi1300m;
wire cdxi1302m = cdxi361m&cdxi445m ^ r83m;
wire cdxi1303m = cdxi405m&cdxi240m;
wire cdxi1304m = cdxi219m&cdxi445m;
wire cdxi1305m = cdxi1303m&r1m;
wire cdxi1306m = cdxi504m&cdxi311m;
wire cdxi1307m = cdxi361m&cdxi241m;
wire cdxi1308m = cdxi361m&cdxi242m;
wire cdxi1309m = cdxi445m&r13m;
wire cdxi1310m = cdxi184m&cdxi528m;
wire cdxi1311m = cdxi405m&r15m;
wire cdxi1312m = cdxi524m&r18m;
wire cdxi1313m = cdxi504m&r19m;
wire cdxi1314m = cdxi361m&r22m;
wire cdxi1315m = cdxi240m&r43m;
wire cdxi1316m = cdxi196m&r44m;
wire cdxi1317m = cdxi184m&r47m;
wire cdxi1318m = cdxi219m&r53m;
wire cdxi1319m = (cdxi1302m ^ cdxi1305m ^ cdxi1306m ^ cdxi1307m ^ cdxi1308m ^ cdxi1309m ^ cdxi1310m ^ cdxi1311m ^ cdxi1312m ^ cdxi1313m ^ cdxi1314m ^ cdxi1315m ^ cdxi1316m ^ cdxi1317m ^ cdxi1318m);
wire cdxi1320m = a0&cdxi1319m;
wire cdxi1321m = (reg_0_91);
wire cdxi1322m = reg_0_3&cdxi535m;
wire cdxi1323m = reg_0_2&cdxi592m;
wire cdxi1324m = reg_0_2&cdxi593m;
wire cdxi1325m = reg_0_2&cdxi594m;
wire cdxi1326m = reg_0_4&cdxi688m;
wire cdxi1327m = reg_0_3&cdxi538m;
wire cdxi1328m = reg_0_3&cdxi539m;
wire cdxi1329m = reg_0_2&cdxi595m;
wire cdxi1330m = reg_0_2&cdxi596m;
wire cdxi1331m = reg_0_2&cdxi597m;
wire cdxi1332m = reg_0_5&cdxi514m;
wire cdxi1333m = reg_0_4&cdxi684m;
wire cdxi1334m = reg_0_3&cdxi534m;
wire cdxi1335m = reg_0_2&cdxi591m;
wire cdxi1336m = (cdxi1322m ^ cdxi1323m ^ cdxi1324m ^ cdxi1325m ^ cdxi1326m ^ cdxi1327m ^ cdxi1328m ^ cdxi1329m ^ cdxi1330m ^ cdxi1331m ^ cdxi1332m ^ cdxi1333m ^ cdxi1334m ^ cdxi1335m ^ cdxi1321m);
wire cdxi1337m = reg_0_0&cdxi1336m;
wire cdxi1338m = cdxi361m&cdxi562m ^ r85m;
wire cdxi1339m = cdxi504m&cdxi207m;
wire cdxi1340m = cdxi405m&cdxi271m;
wire cdxi1341m = cdxi504m&cdxi230m;
wire cdxi1342m = cdxi361m&cdxi325m;
wire cdxi1343m = cdxi361m&cdxi326m;
wire cdxi1344m = cdxi562m&r13m;
wire cdxi1345m = cdxi425m&r14m;
wire cdxi1346m = cdxi405m&r17m;
wire cdxi1347m = cdxi563m&r18m;
wire cdxi1348m = cdxi504m&r21m;
wire cdxi1349m = cdxi361m&r24m;
wire cdxi1350m = cdxi207m&r43m;
wire cdxi1351m = cdxi196m&r46m;
wire cdxi1352m = cdxi184m&r49m;
wire cdxi1353m = cdxi219m&r55m;
wire cdxi1354m = (cdxi1338m ^ cdxi1340m ^ cdxi1341m ^ cdxi1342m ^ cdxi1343m ^ cdxi1344m ^ cdxi1345m ^ cdxi1346m ^ cdxi1347m ^ cdxi1348m ^ cdxi1349m ^ cdxi1350m ^ cdxi1351m ^ cdxi1352m ^ cdxi1353m);
wire cdxi1355m = a0&cdxi1354m;
wire cdxi1356m = (reg_0_93);
wire cdxi1357m = reg_0_3&cdxi573m;
wire cdxi1358m = reg_0_2&cdxi787m;
wire cdxi1359m = reg_0_2&cdxi788m;
wire cdxi1360m = reg_0_2&cdxi789m;
wire cdxi1361m = reg_0_4&reg_0_7&cdxi373m;
wire cdxi1362m = reg_0_3&cdxi576m;
wire cdxi1363m = reg_0_3&cdxi577m;
wire cdxi1364m = reg_0_2&cdxi790m;
wire cdxi1365m = reg_0_2&cdxi791m;
wire cdxi1366m = reg_0_2&cdxi792m;
wire cdxi1367m = reg_0_7&cdxi514m;
wire cdxi1368m = reg_0_4&cdxi958m;
wire cdxi1369m = reg_0_3&cdxi572m;
wire cdxi1370m = reg_0_2&cdxi786m;
wire cdxi1371m = (cdxi1357m ^ cdxi1358m ^ cdxi1359m ^ cdxi1360m ^ cdxi1361m ^ cdxi1362m ^ cdxi1363m ^ cdxi1364m ^ cdxi1365m ^ cdxi1366m ^ cdxi1367m ^ cdxi1368m ^ cdxi1369m ^ cdxi1370m ^ cdxi1356m);
wire cdxi1372m = reg_0_0&cdxi1371m;
wire cdxi1373m = cdxi361m&cdxi638m ^ r86m;
wire cdxi1374m = cdxi582m&cdxi218m;
wire cdxi1375m = cdxi582m&cdxi220m;
wire cdxi1376m = cdxi524m&cdxi291m;
wire cdxi1377m = cdxi361m&cdxi251m;
wire cdxi1378m = cdxi361m&cdxi252m;
wire cdxi1379m = cdxi638m&r13m;
wire cdxi1380m = cdxi601m&r15m;
wire cdxi1381m = cdxi582m&r16m;
wire cdxi1382m = cdxi384m&r19m;
wire cdxi1383m = cdxi524m&r20m;
wire cdxi1384m = cdxi361m&r25m;
wire cdxi1385m = cdxi218m&r44m;
wire cdxi1386m = cdxi240m&r45m;
wire cdxi1387m = cdxi184m&r50m;
wire cdxi1388m = cdxi219m&r56m;
wire cdxi1389m = (cdxi1373m ^ cdxi1375m ^ cdxi1376m ^ cdxi1377m ^ cdxi1378m ^ cdxi1379m ^ cdxi1380m ^ cdxi1381m ^ cdxi1382m ^ cdxi1383m ^ cdxi1384m ^ cdxi1385m ^ cdxi1386m ^ cdxi1387m ^ cdxi1388m);
wire cdxi1390m = a0&cdxi1389m;
wire cdxi1391m = (reg_0_64);
wire cdxi1392m = (reg_0_94);
wire cdxi1393m = reg_0_3&cdxi725m;
wire cdxi1394m = reg_0_2&reg_0_5&cdxi296m;
wire cdxi1395m = reg_0_2&reg_0_3&cdxi256m;
wire cdxi1396m = reg_0_2&reg_0_3&cdxi257m;
wire cdxi1397m = reg_0_5&cdxi706m;
wire cdxi1398m = reg_0_3&cdxi728m;
wire cdxi1399m = reg_0_3&cdxi729m;
wire cdxi1400m = reg_0_2&reg_0_6&cdxi315m;
wire cdxi1401m = reg_0_2&reg_0_5&cdxi295m;
wire cdxi1402m = reg_0_2&reg_0_3&cdxi255m;
wire cdxi1403m = reg_0_6&cdxi684m;
wire cdxi1404m = reg_0_5&cdxi702m;
wire cdxi1405m = reg_0_3&cdxi724m;
wire cdxi1406m = reg_0_2&cdxi1391m;
wire cdxi1407m = (cdxi1393m ^ cdxi1394m ^ cdxi1395m ^ cdxi1396m ^ cdxi1397m ^ cdxi1398m ^ cdxi1399m ^ cdxi1400m ^ cdxi1401m ^ cdxi1402m ^ cdxi1403m ^ cdxi1404m ^ cdxi1405m ^ cdxi1406m ^ cdxi1392m);
wire cdxi1408m = reg_0_0&cdxi1407m;
wire cdxi1409m = cdxi361m&cdxi485m ^ r87m;
wire cdxi1410m = cdxi219m&cdxi485m;
wire cdxi1411m = cdxi582m&cdxi271m;
wire cdxi1412m = cdxi524m&cdxi230m;
wire cdxi1413m = cdxi361m&cdxi261m;
wire cdxi1414m = cdxi361m&cdxi262m;
wire cdxi1415m = cdxi485m&r13m;
wire cdxi1416m = cdxi425m&r15m;
wire cdxi1417m = cdxi582m&r17m;
wire cdxi1418m = cdxi563m&r19m;
wire cdxi1419m = cdxi524m&r21m;
wire cdxi1420m = cdxi361m&r26m;
wire cdxi1421m = cdxi207m&r44m;
wire cdxi1422m = cdxi240m&r46m;
wire cdxi1423m = cdxi184m&r51m;
wire cdxi1424m = cdxi219m&r57m;
wire cdxi1425m = (cdxi1409m ^ cdxi1411m ^ cdxi1412m ^ cdxi1413m ^ cdxi1414m ^ cdxi1415m ^ cdxi1416m ^ cdxi1417m ^ cdxi1418m ^ cdxi1419m ^ cdxi1420m ^ cdxi1421m ^ cdxi1422m ^ cdxi1423m ^ cdxi1424m);
wire cdxi1426m = a0&cdxi1425m;
wire cdxi1427m = (reg_0_95);
wire cdxi1428m = reg_0_3&cdxi743m;
wire cdxi1429m = reg_0_2&cdxi629m;
wire cdxi1430m = reg_0_2&cdxi630m;
wire cdxi1431m = reg_0_2&cdxi631m;
wire cdxi1432m = reg_0_5&reg_0_7&cdxi373m;
wire cdxi1433m = reg_0_3&cdxi746m;
wire cdxi1434m = reg_0_3&cdxi747m;
wire cdxi1435m = reg_0_2&cdxi632m;
wire cdxi1436m = reg_0_2&cdxi633m;
wire cdxi1437m = reg_0_2&cdxi634m;
wire cdxi1438m = reg_0_7&cdxi684m;
wire cdxi1439m = reg_0_5&cdxi958m;
wire cdxi1440m = reg_0_3&cdxi742m;
wire cdxi1441m = reg_0_2&cdxi628m;
wire cdxi1442m = (cdxi1428m ^ cdxi1429m ^ cdxi1430m ^ cdxi1431m ^ cdxi1432m ^ cdxi1433m ^ cdxi1434m ^ cdxi1435m ^ cdxi1436m ^ cdxi1437m ^ cdxi1438m ^ cdxi1439m ^ cdxi1440m ^ cdxi1441m ^ cdxi1427m);
wire cdxi1443m = reg_0_0&cdxi1442m;
wire cdxi1444m = cdxi361m&cdxi657m ^ r88m;
wire cdxi1445m = cdxi601m&cdxi271m;
wire cdxi1446m = cdxi384m&cdxi230m;
wire cdxi1447m = cdxi361m&cdxi337m;
wire cdxi1448m = cdxi361m&cdxi338m;
wire cdxi1449m = cdxi657m&r13m;
wire cdxi1450m = cdxi425m&r16m;
wire cdxi1451m = cdxi601m&r17m;
wire cdxi1452m = cdxi563m&r20m;
wire cdxi1453m = cdxi384m&r21m;
wire cdxi1454m = cdxi361m&r27m;
wire cdxi1455m = cdxi207m&r45m;
wire cdxi1456m = cdxi218m&r46m;
wire cdxi1457m = cdxi184m&r52m;
wire cdxi1458m = cdxi219m&r58m;
wire cdxi1459m = (cdxi1444m ^ cdxi1445m ^ cdxi1446m ^ cdxi1447m ^ cdxi1448m ^ cdxi1449m ^ cdxi1450m ^ cdxi1451m ^ cdxi1452m ^ cdxi1453m ^ cdxi1454m ^ cdxi1455m ^ cdxi1456m ^ cdxi1457m ^ cdxi1458m);
wire cdxi1460m = a0&cdxi1459m;
wire cdxi1461m = (reg_0_96);
wire cdxi1462m = reg_0_3&reg_0_6&cdxi276m;
wire cdxi1463m = reg_0_2&reg_0_6&cdxi235m;
wire cdxi1464m = reg_0_2&reg_0_3&cdxi342m;
wire cdxi1465m = reg_0_2&reg_0_3&cdxi343m;
wire cdxi1466m = reg_0_6&reg_0_7&cdxi373m;
wire cdxi1467m = reg_0_3&reg_0_7&cdxi224m;
wire cdxi1468m = reg_0_3&reg_0_6&cdxi275m;
wire cdxi1469m = reg_0_2&reg_0_7&cdxi295m;
wire cdxi1470m = reg_0_2&reg_0_6&cdxi234m;
wire cdxi1471m = reg_0_2&reg_0_3&cdxi341m;
wire cdxi1472m = reg_0_7&cdxi702m;
wire cdxi1473m = reg_0_6&cdxi958m;
wire cdxi1474m = reg_0_3&cdxi1069m;
wire cdxi1475m = reg_0_2&cdxi1213m;
wire cdxi1476m = (cdxi1462m ^ cdxi1463m ^ cdxi1464m ^ cdxi1465m ^ cdxi1466m ^ cdxi1467m ^ cdxi1468m ^ cdxi1469m ^ cdxi1470m ^ cdxi1471m ^ cdxi1472m ^ cdxi1473m ^ cdxi1474m ^ cdxi1475m ^ cdxi1461m);
wire cdxi1477m = reg_0_0&cdxi1476m;
wire cdxi1478m = cdxi1304m&cdxi218m ^ r89m;
wire cdxi1479m = cdxi445m&cdxi218m;
wire cdxi1480m = cdxi445m&cdxi220m;
wire cdxi1481m = cdxi524m&cdxi301m;
wire cdxi1482m = cdxi504m&cdxi251m;
wire cdxi1483m = cdxi504m&cdxi252m;
wire cdxi1484m = cdxi240m&cdxi547m;
wire cdxi1485m = cdxi466m&r15m;
wire cdxi1486m = cdxi445m&r16m;
wire cdxi1487m = cdxi384m&r22m;
wire cdxi1488m = cdxi524m&r23m;
wire cdxi1489m = cdxi504m&r25m;
wire cdxi1490m = cdxi218m&r47m;
wire cdxi1491m = cdxi240m&r48m;
wire cdxi1492m = cdxi196m&r50m;
wire cdxi1493m = cdxi219m&r59m;
wire cdxi1494m = (cdxi1478m ^ cdxi1480m ^ cdxi1481m ^ cdxi1482m ^ cdxi1483m ^ cdxi1484m ^ cdxi1485m ^ cdxi1486m ^ cdxi1487m ^ cdxi1488m ^ cdxi1489m ^ cdxi1490m ^ cdxi1491m ^ cdxi1492m ^ cdxi1493m);
wire cdxi1495m = a0&cdxi1494m;
wire cdxi1496m = (reg_0_97);
wire cdxi1497m = reg_0_4&cdxi725m;
wire cdxi1498m = reg_0_2&cdxi648m;
wire cdxi1499m = reg_0_2&cdxi649m;
wire cdxi1500m = reg_0_2&cdxi650m;
wire cdxi1501m = reg_0_5&cdxi556m;
wire cdxi1502m = reg_0_4&cdxi728m;
wire cdxi1503m = reg_0_4&cdxi729m;
wire cdxi1504m = reg_0_2&cdxi651m;
wire cdxi1505m = reg_0_2&cdxi652m;
wire cdxi1506m = reg_0_2&cdxi653m;
wire cdxi1507m = reg_0_6&cdxi534m;
wire cdxi1508m = reg_0_5&cdxi552m;
wire cdxi1509m = reg_0_4&cdxi724m;
wire cdxi1510m = reg_0_2&cdxi647m;
wire cdxi1511m = (cdxi1497m ^ cdxi1498m ^ cdxi1499m ^ cdxi1500m ^ cdxi1501m ^ cdxi1502m ^ cdxi1503m ^ cdxi1504m ^ cdxi1505m ^ cdxi1506m ^ cdxi1507m ^ cdxi1508m ^ cdxi1509m ^ cdxi1510m ^ cdxi1496m);
wire cdxi1512m = reg_0_0&cdxi1511m;
wire cdxi1513m = cdxi219m&cdxi1232m ^ r90m;
wire cdxi1514m = cdxi445m&cdxi271m;
wire cdxi1515m = cdxi524m&cdxi325m;
wire cdxi1516m = cdxi504m&cdxi261m;
wire cdxi1517m = cdxi504m&cdxi262m;
wire cdxi1518m = cdxi485m&r14m;
wire cdxi1519m = cdxi562m&r15m;
wire cdxi1520m = cdxi445m&r17m;
wire cdxi1521m = cdxi563m&r22m;
wire cdxi1522m = cdxi524m&r24m;
wire cdxi1523m = cdxi504m&r26m;
wire cdxi1524m = cdxi207m&r47m;
wire cdxi1525m = cdxi240m&r49m;
wire cdxi1526m = cdxi196m&r51m;
wire cdxi1527m = cdxi219m&r60m;
wire cdxi1528m = (cdxi1513m ^ cdxi1514m ^ cdxi1515m ^ cdxi1516m ^ cdxi1517m ^ cdxi1518m ^ cdxi1519m ^ cdxi1520m ^ cdxi1521m ^ cdxi1522m ^ cdxi1523m ^ cdxi1524m ^ cdxi1525m ^ cdxi1526m ^ cdxi1527m);
wire cdxi1529m = a0&cdxi1528m;
wire cdxi1530m = (reg_0_98);
wire cdxi1531m = reg_0_4&cdxi743m;
wire cdxi1532m = reg_0_2&cdxi811m;
wire cdxi1533m = reg_0_2&cdxi812m;
wire cdxi1534m = reg_0_2&cdxi813m;
wire cdxi1535m = reg_0_5&cdxi576m;
wire cdxi1536m = reg_0_4&cdxi746m;
wire cdxi1537m = reg_0_4&cdxi747m;
wire cdxi1538m = reg_0_2&cdxi814m;
wire cdxi1539m = reg_0_2&cdxi815m;
wire cdxi1540m = reg_0_2&cdxi816m;
wire cdxi1541m = reg_0_7&cdxi534m;
wire cdxi1542m = reg_0_5&cdxi572m;
wire cdxi1543m = reg_0_4&cdxi742m;
wire cdxi1544m = reg_0_2&cdxi810m;
wire cdxi1545m = (cdxi1531m ^ cdxi1532m ^ cdxi1533m ^ cdxi1534m ^ cdxi1535m ^ cdxi1536m ^ cdxi1537m ^ cdxi1538m ^ cdxi1539m ^ cdxi1540m ^ cdxi1541m ^ cdxi1542m ^ cdxi1543m ^ cdxi1544m ^ cdxi1530m);
wire cdxi1546m = reg_0_0&cdxi1545m;
wire cdxi1547m = cdxi582m&cdxi657m ^ r96m;
wire cdxi1548m = cdxi638m&cdxi207m;
wire cdxi1549m = cdxi638m&cdxi230m;
wire cdxi1550m = cdxi601m&cdxi261m;
wire cdxi1551m = cdxi582m&cdxi337m;
wire cdxi1552m = cdxi582m&cdxi338m;
wire cdxi1553m = cdxi218m&cdxi623m;
wire cdxi1554m = cdxi485m&r20m;
wire cdxi1555m = cdxi638m&r21m;
wire cdxi1556m = cdxi425m&r25m;
wire cdxi1557m = cdxi601m&r26m;
wire cdxi1558m = cdxi582m&r27m;
wire cdxi1559m = cdxi207m&r56m;
wire cdxi1560m = cdxi218m&r57m;
wire cdxi1561m = cdxi240m&r58m;
wire cdxi1562m = cdxi184m&r62m;
wire cdxi1563m = (cdxi1547m ^ cdxi1549m ^ cdxi1550m ^ cdxi1551m ^ cdxi1552m ^ cdxi1553m ^ cdxi1554m ^ cdxi1555m ^ cdxi1556m ^ cdxi1557m ^ cdxi1558m ^ cdxi1559m ^ cdxi1560m ^ cdxi1561m ^ cdxi1562m);
wire cdxi1564m = a0&cdxi1563m;
wire cdxi1565m = (reg_0_104);
wire cdxi1566m = reg_0_5&reg_0_6&cdxi235m;
wire cdxi1567m = reg_0_3&cdxi667m;
wire cdxi1568m = reg_0_3&cdxi668m;
wire cdxi1569m = reg_0_3&cdxi669m;
wire cdxi1570m = reg_0_6&cdxi632m;
wire cdxi1571m = reg_0_5&reg_0_7&cdxi295m;
wire cdxi1572m = reg_0_5&reg_0_6&cdxi234m;
wire cdxi1573m = reg_0_3&cdxi670m;
wire cdxi1574m = reg_0_3&cdxi671m;
wire cdxi1575m = reg_0_3&cdxi672m;
wire cdxi1576m = reg_0_7&cdxi1391m;
wire cdxi1577m = reg_0_6&cdxi628m;
wire cdxi1578m = reg_0_5&cdxi1213m;
wire cdxi1579m = reg_0_3&cdxi666m;
wire cdxi1580m = (cdxi1566m ^ cdxi1567m ^ cdxi1568m ^ cdxi1569m ^ cdxi1570m ^ cdxi1571m ^ cdxi1572m ^ cdxi1573m ^ cdxi1574m ^ cdxi1575m ^ cdxi1576m ^ cdxi1577m ^ cdxi1578m ^ cdxi1579m ^ cdxi1565m);
wire cdxi1581m = reg_0_0&cdxi1580m;
wire cdxi1582m = cdxi361m&cdxi466m ^ r84m;
wire cdxi1583m = cdxi405m&cdxi220m;
wire cdxi1584m = cdxi504m&cdxi291m;
wire cdxi1585m = cdxi361m&cdxi301m;
wire cdxi1586m = cdxi361m&cdxi302m;
wire cdxi1587m = cdxi466m&r13m;
wire cdxi1588m = cdxi184m&cdxi547m;
wire cdxi1589m = cdxi405m&r16m;
wire cdxi1590m = cdxi384m&r18m;
wire cdxi1591m = cdxi504m&r20m;
wire cdxi1592m = cdxi361m&r23m;
wire cdxi1593m = cdxi218m&r43m;
wire cdxi1594m = cdxi196m&r45m;
wire cdxi1595m = cdxi184m&r48m;
wire cdxi1596m = cdxi219m&r54m;
wire cdxi1597m = (cdxi1582m ^ cdxi1583m ^ cdxi1584m ^ cdxi1585m ^ cdxi1586m ^ cdxi1587m ^ cdxi1588m ^ cdxi1589m ^ cdxi1590m ^ cdxi1591m ^ cdxi1592m ^ cdxi1593m ^ cdxi1594m ^ cdxi1595m ^ cdxi1596m);
wire cdxi1598m = cdxi185m&cdxi1597m;
wire cdxi1599m = (reg_0_92);
wire cdxi1600m = reg_0_3&cdxi553m;
wire cdxi1601m = reg_0_2&cdxi611m;
wire cdxi1602m = reg_0_2&cdxi612m;
wire cdxi1603m = reg_0_2&cdxi613m;
wire cdxi1604m = reg_0_4&cdxi706m;
wire cdxi1605m = reg_0_3&cdxi556m;
wire cdxi1606m = reg_0_3&cdxi557m;
wire cdxi1607m = reg_0_2&cdxi614m;
wire cdxi1608m = reg_0_2&cdxi615m;
wire cdxi1609m = reg_0_2&cdxi616m;
wire cdxi1610m = reg_0_6&cdxi514m;
wire cdxi1611m = reg_0_4&cdxi702m;
wire cdxi1612m = reg_0_3&cdxi552m;
wire cdxi1613m = reg_0_2&cdxi610m;
wire cdxi1614m = (cdxi1600m ^ cdxi1601m ^ cdxi1602m ^ cdxi1603m ^ cdxi1604m ^ cdxi1605m ^ cdxi1606m ^ cdxi1607m ^ cdxi1608m ^ cdxi1609m ^ cdxi1610m ^ cdxi1611m ^ cdxi1612m ^ cdxi1613m ^ cdxi1599m);
wire cdxi1615m = reg_0_1&cdxi1614m;
wire cdxi1616m = cdxi185m&cdxi1528m;
wire cdxi1617m = reg_0_1&cdxi1545m;
wire cdxi1618m = cdxi405m&cdxi485m ^ r94m;
wire cdxi1619m = cdxi445m&cdxi230m;
wire cdxi1620m = cdxi582m&cdxi325m;
wire cdxi1621m = cdxi405m&cdxi261m;
wire cdxi1622m = cdxi405m&cdxi262m;
wire cdxi1623m = cdxi485m&r18m;
wire cdxi1624m = cdxi562m&r19m;
wire cdxi1625m = cdxi445m&r21m;
wire cdxi1626m = cdxi425m&r22m;
wire cdxi1627m = cdxi582m&r24m;
wire cdxi1628m = cdxi405m&r26m;
wire cdxi1629m = cdxi207m&r53m;
wire cdxi1630m = cdxi240m&r55m;
wire cdxi1631m = cdxi196m&r57m;
wire cdxi1632m = cdxi184m&r60m;
wire cdxi1633m = (cdxi1618m ^ cdxi1619m ^ cdxi1620m ^ cdxi1621m ^ cdxi1622m ^ cdxi1623m ^ cdxi1624m ^ cdxi1625m ^ cdxi1626m ^ cdxi1627m ^ cdxi1628m ^ cdxi1629m ^ cdxi1630m ^ cdxi1631m ^ cdxi1632m);
wire cdxi1634m = cdxi185m&cdxi1633m;
wire cdxi1635m = (reg_0_102);
wire cdxi1636m = reg_0_4&cdxi629m;
wire cdxi1637m = reg_0_3&cdxi811m;
wire cdxi1638m = reg_0_3&cdxi812m;
wire cdxi1639m = reg_0_3&cdxi813m;
wire cdxi1640m = reg_0_5&cdxi790m;
wire cdxi1641m = reg_0_4&cdxi632m;
wire cdxi1642m = reg_0_4&cdxi633m;
wire cdxi1643m = reg_0_3&cdxi814m;
wire cdxi1644m = reg_0_3&cdxi815m;
wire cdxi1645m = reg_0_3&cdxi816m;
wire cdxi1646m = reg_0_7&cdxi591m;
wire cdxi1647m = reg_0_5&cdxi786m;
wire cdxi1648m = reg_0_4&cdxi628m;
wire cdxi1649m = reg_0_3&cdxi810m;
wire cdxi1650m = (cdxi1636m ^ cdxi1637m ^ cdxi1638m ^ cdxi1639m ^ cdxi1640m ^ cdxi1641m ^ cdxi1642m ^ cdxi1643m ^ cdxi1644m ^ cdxi1645m ^ cdxi1646m ^ cdxi1647m ^ cdxi1648m ^ cdxi1649m ^ cdxi1635m);
wire cdxi1651m = reg_0_1&cdxi1650m;
wire cdxi1652m = cdxi405m&cdxi657m ^ r95m;
wire cdxi1653m = cdxi466m&cdxi230m;
wire cdxi1654m = cdxi601m&cdxi325m;
wire cdxi1655m = cdxi405m&cdxi337m;
wire cdxi1656m = cdxi405m&cdxi338m;
wire cdxi1657m = cdxi657m&r18m;
wire cdxi1658m = cdxi562m&r20m;
wire cdxi1659m = cdxi466m&r21m;
wire cdxi1660m = cdxi425m&r23m;
wire cdxi1661m = cdxi601m&r24m;
wire cdxi1662m = cdxi405m&r27m;
wire cdxi1663m = cdxi207m&r54m;
wire cdxi1664m = cdxi218m&r55m;
wire cdxi1665m = cdxi196m&r58m;
wire cdxi1666m = cdxi184m&r61m;
wire cdxi1667m = (cdxi1652m ^ cdxi1653m ^ cdxi1654m ^ cdxi1655m ^ cdxi1656m ^ cdxi1657m ^ cdxi1658m ^ cdxi1659m ^ cdxi1660m ^ cdxi1661m ^ cdxi1662m ^ cdxi1663m ^ cdxi1664m ^ cdxi1665m ^ cdxi1666m);
wire cdxi1668m = cdxi185m&cdxi1667m;
wire cdxi1669m = (reg_0_103);
wire cdxi1670m = reg_0_4&reg_0_6&cdxi235m;
wire cdxi1671m = reg_0_3&cdxi767m;
wire cdxi1672m = reg_0_3&cdxi768m;
wire cdxi1673m = reg_0_3&cdxi769m;
wire cdxi1674m = reg_0_6&cdxi790m;
wire cdxi1675m = reg_0_4&reg_0_7&cdxi295m;
wire cdxi1676m = reg_0_4&reg_0_6&cdxi234m;
wire cdxi1677m = reg_0_3&cdxi770m;
wire cdxi1678m = reg_0_3&cdxi771m;
wire cdxi1679m = reg_0_3&cdxi772m;
wire cdxi1680m = reg_0_7&cdxi610m;
wire cdxi1681m = reg_0_6&cdxi786m;
wire cdxi1682m = reg_0_4&cdxi1213m;
wire cdxi1683m = reg_0_3&cdxi766m;
wire cdxi1684m = (cdxi1670m ^ cdxi1671m ^ cdxi1672m ^ cdxi1673m ^ cdxi1674m ^ cdxi1675m ^ cdxi1676m ^ cdxi1677m ^ cdxi1678m ^ cdxi1679m ^ cdxi1680m ^ cdxi1681m ^ cdxi1682m ^ cdxi1683m ^ cdxi1669m);
wire cdxi1685m = reg_0_1&cdxi1684m;
wire cdxi1686m = cdxi405m&cdxi638m ^ r93m;
wire cdxi1687m = cdxi445m&cdxi291m;
wire cdxi1688m = cdxi582m&cdxi301m;
wire cdxi1689m = cdxi405m&cdxi251m;
wire cdxi1690m = cdxi405m&cdxi252m;
wire cdxi1691m = cdxi240m&cdxi605m;
wire cdxi1692m = cdxi466m&r19m;
wire cdxi1693m = cdxi445m&r20m;
wire cdxi1694m = cdxi601m&r22m;
wire cdxi1695m = cdxi582m&r23m;
wire cdxi1696m = cdxi405m&r25m;
wire cdxi1697m = cdxi218m&r53m;
wire cdxi1698m = cdxi240m&r54m;
wire cdxi1699m = cdxi196m&r56m;
wire cdxi1700m = cdxi184m&r59m;
wire cdxi1701m = (cdxi1686m ^ cdxi1687m ^ cdxi1688m ^ cdxi1689m ^ cdxi1690m ^ cdxi1691m ^ cdxi1692m ^ cdxi1693m ^ cdxi1694m ^ cdxi1695m ^ cdxi1696m ^ cdxi1697m ^ cdxi1698m ^ cdxi1699m ^ cdxi1700m);
wire cdxi1702m = cdxi219m&cdxi1701m;
wire cdxi1703m = (reg_0_101);
wire cdxi1704m = reg_0_4&reg_0_5&cdxi296m;
wire cdxi1705m = reg_0_3&cdxi648m;
wire cdxi1706m = reg_0_3&cdxi649m;
wire cdxi1707m = reg_0_3&cdxi650m;
wire cdxi1708m = reg_0_5&cdxi614m;
wire cdxi1709m = reg_0_4&reg_0_6&cdxi315m;
wire cdxi1710m = reg_0_4&reg_0_5&cdxi295m;
wire cdxi1711m = reg_0_3&cdxi651m;
wire cdxi1712m = reg_0_3&cdxi652m;
wire cdxi1713m = reg_0_3&cdxi653m;
wire cdxi1714m = reg_0_6&cdxi591m;
wire cdxi1715m = reg_0_5&cdxi610m;
wire cdxi1716m = reg_0_4&cdxi1391m;
wire cdxi1717m = reg_0_3&cdxi647m;
wire cdxi1718m = (cdxi1704m ^ cdxi1705m ^ cdxi1706m ^ cdxi1707m ^ cdxi1708m ^ cdxi1709m ^ cdxi1710m ^ cdxi1711m ^ cdxi1712m ^ cdxi1713m ^ cdxi1714m ^ cdxi1715m ^ cdxi1716m ^ cdxi1717m ^ cdxi1703m);
wire cdxi1719m = reg_0_2&cdxi1718m;
wire cdxi1720m = cdxi219m&cdxi1633m;
wire cdxi1721m = reg_0_2&cdxi1650m;
wire cdxi1722m = cdxi219m&cdxi1667m;
wire cdxi1723m = reg_0_2&cdxi1684m;
wire cdxi1724m = cdxi219m&cdxi1563m;
wire cdxi1725m = reg_0_2&cdxi1580m;
wire cdxi1726m = cdxi445m&cdxi657m ^ r97m;
wire cdxi1727m = cdxi638m&cdxi325m;
wire cdxi1728m = cdxi466m&cdxi261m;
wire cdxi1729m = cdxi445m&cdxi337m;
wire cdxi1730m = cdxi445m&cdxi338m;
wire cdxi1731m = cdxi657m&r22m;
wire cdxi1732m = cdxi485m&r23m;
wire cdxi1733m = cdxi638m&r24m;
wire cdxi1734m = cdxi562m&r25m;
wire cdxi1735m = cdxi466m&r26m;
wire cdxi1736m = cdxi445m&r27m;
wire cdxi1737m = cdxi207m&r59m;
wire cdxi1738m = cdxi218m&r60m;
wire cdxi1739m = cdxi240m&r61m;
wire cdxi1740m = cdxi196m&r62m;
wire cdxi1741m = (cdxi1726m ^ cdxi1727m ^ cdxi1728m ^ cdxi1729m ^ cdxi1730m ^ cdxi1731m ^ cdxi1732m ^ cdxi1733m ^ cdxi1734m ^ cdxi1735m ^ cdxi1736m ^ cdxi1737m ^ cdxi1738m ^ cdxi1739m ^ cdxi1740m);
wire cdxi1742m = cdxi184m&cdxi1741m;
wire cdxi1743m = (reg_0_105);
wire cdxi1744m = reg_0_5&cdxi767m;
wire cdxi1745m = reg_0_4&cdxi667m;
wire cdxi1746m = reg_0_4&cdxi668m;
wire cdxi1747m = reg_0_4&cdxi669m;
wire cdxi1748m = reg_0_6&cdxi814m;
wire cdxi1749m = reg_0_5&cdxi770m;
wire cdxi1750m = reg_0_5&cdxi771m;
wire cdxi1751m = reg_0_4&cdxi670m;
wire cdxi1752m = reg_0_4&cdxi671m;
wire cdxi1753m = reg_0_4&cdxi672m;
wire cdxi1754m = reg_0_7&cdxi647m;
wire cdxi1755m = reg_0_6&cdxi810m;
wire cdxi1756m = reg_0_5&cdxi766m;
wire cdxi1757m = reg_0_4&cdxi666m;
wire cdxi1758m = (cdxi1744m ^ cdxi1745m ^ cdxi1746m ^ cdxi1747m ^ cdxi1748m ^ cdxi1749m ^ cdxi1750m ^ cdxi1751m ^ cdxi1752m ^ cdxi1753m ^ cdxi1754m ^ cdxi1755m ^ cdxi1756m ^ cdxi1757m ^ cdxi1743m);
wire cdxi1759m = reg_0_3&cdxi1758m;
wire cdxi1760m = cdxi825m&cdxi445m ^ r98m;
wire cdxi1761m = cdxi361m&cdxi445m;
wire cdxi1762m = cdxi362m&cdxi445m;
wire cdxi1763m = cdxi363m&cdxi445m;
wire cdxi1764m = cdxi825m&cdxi240m;
wire cdxi1765m = cdxi185m&cdxi822m;
wire cdxi1766m = cdxi361m&cdxi447m;
wire cdxi1767m = cdxi362m&cdxi525m;
wire cdxi1768m = cdxi363m&cdxi583m;
wire cdxi1769m = cdxi825m&cdxi241m;
wire cdxi1770m = cdxi825m&cdxi242m;
wire cdxi1771m = cdxi1303m&r7m;
wire cdxi1772m = cdxi1304m&r8m;
wire cdxi1773m = cdxi361m&cdxi450m;
wire cdxi1774m = cdxi361m&cdxi451m;
wire cdxi1775m = cdxi406m&cdxi679m;
wire cdxi1776m = cdxi362m&cdxi528m;
wire cdxi1777m = cdxi362m&cdxi529m;
wire cdxi1778m = cdxi363m&cdxi586m;
wire cdxi1779m = cdxi363m&cdxi587m;
wire cdxi1780m = cdxi825m&r22m;
wire cdxi1781m = cdxi445m&r28m;
wire cdxi1782m = cdxi582m&r29m;
wire cdxi1783m = cdxi405m&r30m;
wire cdxi1784m = cdxi524m&r33m;
wire cdxi1785m = cdxi504m&r34m;
wire cdxi1786m = cdxi361m&r37m;
wire cdxi1787m = cdxi446m&r43m;
wire cdxi1788m = cdxi406m&r44m;
wire cdxi1789m = cdxi362m&r47m;
wire cdxi1790m = cdxi363m&r53m;
wire cdxi1791m = cdxi240m&r63m;
wire cdxi1792m = cdxi196m&r64m;
wire cdxi1793m = cdxi184m&r67m;
wire cdxi1794m = cdxi219m&r73m;
wire cdxi1795m = cdxi185m&r83m;
wire cdxi1796m = (cdxi1760m ^ cdxi1766m ^ cdxi1767m ^ cdxi1768m ^ cdxi1769m ^ cdxi1770m ^ cdxi1771m ^ cdxi1772m ^ cdxi1773m ^ cdxi1774m ^ cdxi1775m ^ cdxi1776m ^ cdxi1777m ^ cdxi1778m ^ cdxi1779m ^ cdxi1780m ^ cdxi1781m ^ cdxi1782m ^ cdxi1783m ^ cdxi1784m ^ cdxi1785m ^ cdxi1786m ^ cdxi1787m ^ cdxi1788m ^ cdxi1789m ^ cdxi1790m ^ cdxi1791m ^ cdxi1792m ^ cdxi1793m ^ cdxi1794m ^ cdxi1795m);
wire cdxi1797m = a0&cdxi1796m;
wire cdxi1798m = (reg_0_75);
wire cdxi1799m = (reg_0_81);
wire cdxi1800m = (reg_0_106);
wire cdxi1801m = reg_0_2&reg_0_3&cdxi457m;
wire cdxi1802m = reg_0_1&cdxi1322m;
wire cdxi1803m = reg_0_1&cdxi1323m;
wire cdxi1804m = reg_0_1&cdxi1324m;
wire cdxi1805m = reg_0_1&cdxi1325m;
wire cdxi1806m = reg_0_3&reg_0_4&reg_0_5&cdxi372m;
wire cdxi1807m = reg_0_2&reg_0_4&reg_0_5&cdxi190m;
wire cdxi1808m = reg_0_2&reg_0_3&cdxi460m;
wire cdxi1809m = reg_0_2&reg_0_3&cdxi461m;
wire cdxi1810m = reg_0_1&cdxi1326m;
wire cdxi1811m = reg_0_1&cdxi1327m;
wire cdxi1812m = reg_0_1&cdxi1328m;
wire cdxi1813m = reg_0_1&cdxi1329m;
wire cdxi1814m = reg_0_1&cdxi1330m;
wire cdxi1815m = reg_0_1&cdxi1331m;
wire cdxi1816m = reg_0_4&cdxi893m;
wire cdxi1817m = reg_0_3&reg_0_5&cdxi842m;
wire cdxi1818m = reg_0_3&reg_0_4&cdxi880m;
wire cdxi1819m = reg_0_2&reg_0_5&cdxi415m;
wire cdxi1820m = reg_0_2&reg_0_4&cdxi881m;
wire cdxi1821m = reg_0_2&reg_0_3&cdxi456m;
wire cdxi1822m = reg_0_1&cdxi1332m;
wire cdxi1823m = reg_0_1&cdxi1333m;
wire cdxi1824m = reg_0_1&cdxi1334m;
wire cdxi1825m = reg_0_1&cdxi1335m;
wire cdxi1826m = reg_0_5&cdxi843m;
wire cdxi1827m = reg_0_4&cdxi882m;
wire cdxi1828m = reg_0_3&cdxi1798m;
wire cdxi1829m = reg_0_2&cdxi1799m;
wire cdxi1830m = reg_0_1&cdxi1321m;
wire cdxi1831m = (cdxi1801m ^ cdxi1802m ^ cdxi1803m ^ cdxi1804m ^ cdxi1805m ^ cdxi1806m ^ cdxi1807m ^ cdxi1808m ^ cdxi1809m ^ cdxi1810m ^ cdxi1811m ^ cdxi1812m ^ cdxi1813m ^ cdxi1814m ^ cdxi1815m ^ cdxi1816m ^ cdxi1817m ^ cdxi1818m ^ cdxi1819m ^ cdxi1820m ^ cdxi1821m ^ cdxi1822m ^ cdxi1823m ^ cdxi1824m ^ cdxi1825m ^ cdxi1826m ^ cdxi1827m ^ cdxi1828m ^ cdxi1829m ^ cdxi1830m ^ cdxi1800m);
wire cdxi1832m = reg_0_0&cdxi1831m;
wire cdxi1833m = cdxi825m&cdxi466m ^ r99m;
wire cdxi1834m = cdxi361m&cdxi466m;
wire cdxi1835m = cdxi362m&cdxi466m;
wire cdxi1836m = cdxi363m&cdxi466m;
wire cdxi1837m = cdxi825m&cdxi218m;
wire cdxi1838m = cdxi361m&cdxi467m;
wire cdxi1839m = cdxi362m&cdxi544m;
wire cdxi1840m = cdxi363m&cdxi602m;
wire cdxi1841m = cdxi825m&cdxi301m;
wire cdxi1842m = cdxi825m&cdxi302m;
wire cdxi1843m = cdxi405m&cdxi389m;
wire cdxi1844m = cdxi977m&r8m;
wire cdxi1845m = cdxi361m&cdxi470m;
wire cdxi1846m = cdxi361m&cdxi471m;
wire cdxi1847m = cdxi406m&cdxi697m;
wire cdxi1848m = cdxi362m&cdxi547m;
wire cdxi1849m = cdxi362m&cdxi548m;
wire cdxi1850m = cdxi363m&cdxi605m;
wire cdxi1851m = cdxi363m&cdxi606m;
wire cdxi1852m = cdxi825m&r23m;
wire cdxi1853m = cdxi466m&r28m;
wire cdxi1854m = cdxi601m&r29m;
wire cdxi1855m = cdxi405m&r31m;
wire cdxi1856m = cdxi384m&r33m;
wire cdxi1857m = cdxi504m&r35m;
wire cdxi1858m = cdxi361m&r38m;
wire cdxi1859m = cdxi385m&r43m;
wire cdxi1860m = cdxi406m&r45m;
wire cdxi1861m = cdxi362m&r48m;
wire cdxi1862m = cdxi363m&r54m;
wire cdxi1863m = cdxi218m&r63m;
wire cdxi1864m = cdxi196m&r65m;
wire cdxi1865m = cdxi184m&r68m;
wire cdxi1866m = cdxi219m&r74m;
wire cdxi1867m = cdxi185m&r84m;
wire cdxi1868m = (cdxi1833m ^ cdxi1838m ^ cdxi1839m ^ cdxi1840m ^ cdxi1841m ^ cdxi1842m ^ cdxi1843m ^ cdxi1844m ^ cdxi1845m ^ cdxi1846m ^ cdxi1847m ^ cdxi1848m ^ cdxi1849m ^ cdxi1850m ^ cdxi1851m ^ cdxi1852m ^ cdxi1853m ^ cdxi1854m ^ cdxi1855m ^ cdxi1856m ^ cdxi1857m ^ cdxi1858m ^ cdxi1859m ^ cdxi1860m ^ cdxi1861m ^ cdxi1862m ^ cdxi1863m ^ cdxi1864m ^ cdxi1865m ^ cdxi1866m ^ cdxi1867m);
wire cdxi1869m = a0&cdxi1868m;
wire cdxi1870m = (reg_0_107);
wire cdxi1871m = reg_0_2&cdxi1106m;
wire cdxi1872m = reg_0_1&cdxi1600m;
wire cdxi1873m = reg_0_1&cdxi1601m;
wire cdxi1874m = reg_0_1&cdxi1602m;
wire cdxi1875m = reg_0_1&cdxi1603m;
wire cdxi1876m = reg_0_3&cdxi1000m;
wire cdxi1877m = reg_0_2&cdxi1110m;
wire cdxi1878m = reg_0_2&cdxi1111m;
wire cdxi1879m = reg_0_2&cdxi1112m;
wire cdxi1880m = reg_0_1&cdxi1604m;
wire cdxi1881m = reg_0_1&cdxi1605m;
wire cdxi1882m = reg_0_1&cdxi1606m;
wire cdxi1883m = reg_0_1&cdxi1607m;
wire cdxi1884m = reg_0_1&cdxi1608m;
wire cdxi1885m = reg_0_1&cdxi1609m;
wire cdxi1886m = reg_0_4&cdxi931m;
wire cdxi1887m = reg_0_3&cdxi1006m;
wire cdxi1888m = reg_0_3&cdxi1007m;
wire cdxi1889m = reg_0_2&cdxi1116m;
wire cdxi1890m = reg_0_2&cdxi1117m;
wire cdxi1891m = reg_0_2&cdxi1118m;
wire cdxi1892m = reg_0_1&cdxi1610m;
wire cdxi1893m = reg_0_1&cdxi1611m;
wire cdxi1894m = reg_0_1&cdxi1612m;
wire cdxi1895m = reg_0_1&cdxi1613m;
wire cdxi1896m = reg_0_6&cdxi843m;
wire cdxi1897m = reg_0_4&cdxi920m;
wire cdxi1898m = reg_0_3&cdxi995m;
wire cdxi1899m = reg_0_2&cdxi1105m;
wire cdxi1900m = reg_0_1&cdxi1599m;
wire cdxi1901m = (cdxi1871m ^ cdxi1872m ^ cdxi1873m ^ cdxi1874m ^ cdxi1875m ^ cdxi1876m ^ cdxi1877m ^ cdxi1878m ^ cdxi1879m ^ cdxi1880m ^ cdxi1881m ^ cdxi1882m ^ cdxi1883m ^ cdxi1884m ^ cdxi1885m ^ cdxi1886m ^ cdxi1887m ^ cdxi1888m ^ cdxi1889m ^ cdxi1890m ^ cdxi1891m ^ cdxi1892m ^ cdxi1893m ^ cdxi1894m ^ cdxi1895m ^ cdxi1896m ^ cdxi1897m ^ cdxi1898m ^ cdxi1899m ^ cdxi1900m ^ cdxi1870m);
wire cdxi1902m = reg_0_0&cdxi1901m;
wire cdxi1903m = cdxi825m&cdxi638m ^ r101m;
wire cdxi1904m = cdxi361m&cdxi638m;
wire cdxi1905m = cdxi362m&cdxi638m;
wire cdxi1906m = cdxi363m&cdxi638m;
wire cdxi1907m = cdxi1904m&r0m;
wire cdxi1908m = cdxi362m&cdxi716m;
wire cdxi1909m = cdxi863m&cdxi291m;
wire cdxi1910m = cdxi825m&cdxi251m;
wire cdxi1911m = cdxi825m&cdxi252m;
wire cdxi1912m = cdxi582m&cdxi389m;
wire cdxi1913m = cdxi1013m&r8m;
wire cdxi1914m = cdxi900m&r10m;
wire cdxi1915m = cdxi861m&r11m;
wire cdxi1916m = cdxi446m&cdxi697m;
wire cdxi1917m = cdxi362m&cdxi719m;
wire cdxi1918m = cdxi362m&cdxi720m;
wire cdxi1919m = cdxi902m&r19m;
wire cdxi1920m = cdxi863m&r20m;
wire cdxi1921m = cdxi825m&r25m;
wire cdxi1922m = cdxi638m&r28m;
wire cdxi1923m = cdxi601m&r30m;
wire cdxi1924m = cdxi582m&r31m;
wire cdxi1925m = cdxi384m&r34m;
wire cdxi1926m = cdxi524m&r35m;
wire cdxi1927m = cdxi361m&r40m;
wire cdxi1928m = cdxi385m&r44m;
wire cdxi1929m = cdxi446m&r45m;
wire cdxi1930m = cdxi362m&r50m;
wire cdxi1931m = cdxi363m&r56m;
wire cdxi1932m = cdxi218m&r64m;
wire cdxi1933m = cdxi240m&r65m;
wire cdxi1934m = cdxi184m&r70m;
wire cdxi1935m = cdxi219m&r76m;
wire cdxi1936m = cdxi185m&r86m;
wire cdxi1937m = (cdxi1903m ^ cdxi1907m ^ cdxi1908m ^ cdxi1909m ^ cdxi1910m ^ cdxi1911m ^ cdxi1912m ^ cdxi1913m ^ cdxi1914m ^ cdxi1915m ^ cdxi1916m ^ cdxi1917m ^ cdxi1918m ^ cdxi1919m ^ cdxi1920m ^ cdxi1921m ^ cdxi1922m ^ cdxi1923m ^ cdxi1924m ^ cdxi1925m ^ cdxi1926m ^ cdxi1927m ^ cdxi1928m ^ cdxi1929m ^ cdxi1930m ^ cdxi1931m ^ cdxi1932m ^ cdxi1933m ^ cdxi1934m ^ cdxi1935m ^ cdxi1936m);
wire cdxi1938m = a0&cdxi1937m;
wire cdxi1939m = (reg_0_84);
wire cdxi1940m = (reg_0_109);
wire cdxi1941m = reg_0_2&reg_0_3&reg_0_5&reg_0_6&cdxi130m;
wire cdxi1942m = reg_0_1&cdxi1393m;
wire cdxi1943m = reg_0_1&cdxi1394m;
wire cdxi1944m = reg_0_1&cdxi1395m;
wire cdxi1945m = reg_0_1&cdxi1396m;
wire cdxi1946m = reg_0_3&cdxi1037m;
wire cdxi1947m = reg_0_2&reg_0_5&reg_0_6&cdxi190m;
wire cdxi1948m = reg_0_2&reg_0_3&reg_0_6&cdxi455m;
wire cdxi1949m = reg_0_2&reg_0_3&reg_0_5&cdxi394m;
wire cdxi1950m = reg_0_1&cdxi1397m;
wire cdxi1951m = reg_0_1&cdxi1398m;
wire cdxi1952m = reg_0_1&cdxi1399m;
wire cdxi1953m = reg_0_1&cdxi1400m;
wire cdxi1954m = reg_0_1&cdxi1401m;
wire cdxi1955m = reg_0_1&cdxi1402m;
wire cdxi1956m = reg_0_5&cdxi931m;
wire cdxi1957m = reg_0_3&cdxi1043m;
wire cdxi1958m = reg_0_3&cdxi1044m;
wire cdxi1959m = reg_0_2&reg_0_6&cdxi881m;
wire cdxi1960m = reg_0_2&reg_0_5&cdxi919m;
wire cdxi1961m = reg_0_2&reg_0_3&cdxi1031m;
wire cdxi1962m = reg_0_1&cdxi1403m;
wire cdxi1963m = reg_0_1&cdxi1404m;
wire cdxi1964m = reg_0_1&cdxi1405m;
wire cdxi1965m = reg_0_1&cdxi1406m;
wire cdxi1966m = reg_0_6&cdxi882m;
wire cdxi1967m = reg_0_5&cdxi920m;
wire cdxi1968m = reg_0_3&cdxi1032m;
wire cdxi1969m = reg_0_2&cdxi1939m;
wire cdxi1970m = reg_0_1&cdxi1392m;
wire cdxi1971m = (cdxi1941m ^ cdxi1942m ^ cdxi1943m ^ cdxi1944m ^ cdxi1945m ^ cdxi1946m ^ cdxi1947m ^ cdxi1948m ^ cdxi1949m ^ cdxi1950m ^ cdxi1951m ^ cdxi1952m ^ cdxi1953m ^ cdxi1954m ^ cdxi1955m ^ cdxi1956m ^ cdxi1957m ^ cdxi1958m ^ cdxi1959m ^ cdxi1960m ^ cdxi1961m ^ cdxi1962m ^ cdxi1963m ^ cdxi1964m ^ cdxi1965m ^ cdxi1966m ^ cdxi1967m ^ cdxi1968m ^ cdxi1969m ^ cdxi1970m ^ cdxi1940m);
wire cdxi1972m = reg_0_0&cdxi1971m;
wire cdxi1973m = cdxi825m&cdxi485m ^ r102m;
wire cdxi1974m = cdxi361m&cdxi485m;
wire cdxi1975m = cdxi362m&cdxi485m;
wire cdxi1976m = cdxi363m&cdxi485m;
wire cdxi1977m = cdxi825m&cdxi207m;
wire cdxi1978m = cdxi361m&cdxi486m;
wire cdxi1979m = cdxi362m&cdxi734m;
wire cdxi1980m = cdxi363m&cdxi620m;
wire cdxi1981m = cdxi825m&cdxi261m;
wire cdxi1982m = cdxi825m&cdxi262m;
wire cdxi1983m = cdxi1160m&r7m;
wire cdxi1984m = cdxi524m&cdxi430m;
wire cdxi1985m = cdxi361m&cdxi489m;
wire cdxi1986m = cdxi361m&cdxi490m;
wire cdxi1987m = cdxi1161m&r13m;
wire cdxi1988m = cdxi362m&cdxi737m;
wire cdxi1989m = cdxi362m&cdxi738m;
wire cdxi1990m = cdxi363m&cdxi623m;
wire cdxi1991m = cdxi363m&cdxi624m;
wire cdxi1992m = cdxi825m&r26m;
wire cdxi1993m = cdxi485m&r28m;
wire cdxi1994m = cdxi425m&r30m;
wire cdxi1995m = cdxi582m&r32m;
wire cdxi1996m = cdxi563m&r34m;
wire cdxi1997m = cdxi524m&r36m;
wire cdxi1998m = cdxi361m&r41m;
wire cdxi1999m = cdxi426m&r44m;
wire cdxi2000m = cdxi446m&r46m;
wire cdxi2001m = cdxi362m&r51m;
wire cdxi2002m = cdxi363m&r57m;
wire cdxi2003m = cdxi207m&r64m;
wire cdxi2004m = cdxi240m&r66m;
wire cdxi2005m = cdxi184m&r71m;
wire cdxi2006m = cdxi219m&r77m;
wire cdxi2007m = cdxi185m&r87m;
wire cdxi2008m = (cdxi1973m ^ cdxi1978m ^ cdxi1979m ^ cdxi1980m ^ cdxi1981m ^ cdxi1982m ^ cdxi1983m ^ cdxi1984m ^ cdxi1985m ^ cdxi1986m ^ cdxi1987m ^ cdxi1988m ^ cdxi1989m ^ cdxi1990m ^ cdxi1991m ^ cdxi1992m ^ cdxi1993m ^ cdxi1994m ^ cdxi1995m ^ cdxi1996m ^ cdxi1997m ^ cdxi1998m ^ cdxi1999m ^ cdxi2000m ^ cdxi2001m ^ cdxi2002m ^ cdxi2003m ^ cdxi2004m ^ cdxi2005m ^ cdxi2006m ^ cdxi2007m);
wire cdxi2009m = a0&cdxi2008m;
wire cdxi2010m = (reg_0_79);
wire cdxi2011m = (reg_0_110);
wire cdxi2012m = reg_0_2&cdxi1179m;
wire cdxi2013m = reg_0_1&cdxi1428m;
wire cdxi2014m = reg_0_1&cdxi1429m;
wire cdxi2015m = reg_0_1&cdxi1430m;
wire cdxi2016m = reg_0_1&cdxi1431m;
wire cdxi2017m = reg_0_3&reg_0_5&reg_0_7&cdxi372m;
wire cdxi2018m = reg_0_2&cdxi1183m;
wire cdxi2019m = reg_0_2&cdxi1184m;
wire cdxi2020m = reg_0_2&cdxi1185m;
wire cdxi2021m = reg_0_1&cdxi1432m;
wire cdxi2022m = reg_0_1&cdxi1433m;
wire cdxi2023m = reg_0_1&cdxi1434m;
wire cdxi2024m = reg_0_1&cdxi1435m;
wire cdxi2025m = reg_0_1&cdxi1436m;
wire cdxi2026m = reg_0_1&cdxi1437m;
wire cdxi2027m = reg_0_5&cdxi970m;
wire cdxi2028m = reg_0_3&reg_0_7&cdxi880m;
wire cdxi2029m = reg_0_3&reg_0_5&cdxi957m;
wire cdxi2030m = reg_0_2&cdxi1189m;
wire cdxi2031m = reg_0_2&cdxi1190m;
wire cdxi2032m = reg_0_2&cdxi1191m;
wire cdxi2033m = reg_0_1&cdxi1438m;
wire cdxi2034m = reg_0_1&cdxi1439m;
wire cdxi2035m = reg_0_1&cdxi1440m;
wire cdxi2036m = reg_0_1&cdxi1441m;
wire cdxi2037m = reg_0_7&cdxi882m;
wire cdxi2038m = reg_0_5&cdxi959m;
wire cdxi2039m = reg_0_3&cdxi2010m;
wire cdxi2040m = reg_0_2&cdxi1178m;
wire cdxi2041m = reg_0_1&cdxi1427m;
wire cdxi2042m = (cdxi2012m ^ cdxi2013m ^ cdxi2014m ^ cdxi2015m ^ cdxi2016m ^ cdxi2017m ^ cdxi2018m ^ cdxi2019m ^ cdxi2020m ^ cdxi2021m ^ cdxi2022m ^ cdxi2023m ^ cdxi2024m ^ cdxi2025m ^ cdxi2026m ^ cdxi2027m ^ cdxi2028m ^ cdxi2029m ^ cdxi2030m ^ cdxi2031m ^ cdxi2032m ^ cdxi2033m ^ cdxi2034m ^ cdxi2035m ^ cdxi2036m ^ cdxi2037m ^ cdxi2038m ^ cdxi2039m ^ cdxi2040m ^ cdxi2041m ^ cdxi2011m);
wire cdxi2043m = reg_0_0&cdxi2042m;
wire cdxi2044m = cdxi363m&cdxi1479m ^ r104m;
wire cdxi2045m = cdxi1304m&cdxi218m;
wire cdxi2046m = cdxi406m&cdxi638m;
wire cdxi2047m = cdxi2045m&r0m;
wire cdxi2048m = cdxi406m&cdxi716m;
wire cdxi2049m = cdxi363m&cdxi639m;
wire cdxi2050m = cdxi363m&cdxi640m;
wire cdxi2051m = cdxi363m&cdxi641m;
wire cdxi2052m = cdxi445m&cdxi389m;
wire cdxi2053m = cdxi524m&cdxi470m;
wire cdxi2054m = cdxi977m&r10m;
wire cdxi2055m = cdxi1304m&r11m;
wire cdxi2056m = cdxi446m&cdxi547m;
wire cdxi2057m = cdxi406m&cdxi719m;
wire cdxi2058m = cdxi406m&cdxi720m;
wire cdxi2059m = cdxi363m&cdxi642m;
wire cdxi2060m = cdxi363m&cdxi643m;
wire cdxi2061m = cdxi363m&cdxi644m;
wire cdxi2062m = cdxi638m&r29m;
wire cdxi2063m = cdxi466m&r30m;
wire cdxi2064m = cdxi445m&r31m;
wire cdxi2065m = cdxi384m&r37m;
wire cdxi2066m = cdxi524m&r38m;
wire cdxi2067m = cdxi504m&r40m;
wire cdxi2068m = cdxi385m&r47m;
wire cdxi2069m = cdxi446m&r48m;
wire cdxi2070m = cdxi406m&r50m;
wire cdxi2071m = cdxi363m&r59m;
wire cdxi2072m = cdxi218m&r67m;
wire cdxi2073m = cdxi240m&r68m;
wire cdxi2074m = cdxi196m&r70m;
wire cdxi2075m = cdxi219m&r79m;
wire cdxi2076m = cdxi185m&r89m;
wire cdxi2077m = (cdxi2044m ^ cdxi2047m ^ cdxi2048m ^ cdxi2049m ^ cdxi2050m ^ cdxi2051m ^ cdxi2052m ^ cdxi2053m ^ cdxi2054m ^ cdxi2055m ^ cdxi2056m ^ cdxi2057m ^ cdxi2058m ^ cdxi2059m ^ cdxi2060m ^ cdxi2061m ^ cdxi2062m ^ cdxi2063m ^ cdxi2064m ^ cdxi2065m ^ cdxi2066m ^ cdxi2067m ^ cdxi2068m ^ cdxi2069m ^ cdxi2070m ^ cdxi2071m ^ cdxi2072m ^ cdxi2073m ^ cdxi2074m ^ cdxi2075m ^ cdxi2076m);
wire cdxi2078m = a0&cdxi2077m;
wire cdxi2079m = (reg_0_87);
wire cdxi2080m = (reg_0_112);
wire cdxi2081m = reg_0_2&reg_0_4&reg_0_5&reg_0_6&cdxi130m;
wire cdxi2082m = reg_0_1&cdxi1497m;
wire cdxi2083m = reg_0_1&cdxi1498m;
wire cdxi2084m = reg_0_1&cdxi1499m;
wire cdxi2085m = reg_0_1&cdxi1500m;
wire cdxi2086m = reg_0_4&cdxi1037m;
wire cdxi2087m = reg_0_2&reg_0_5&cdxi479m;
wire cdxi2088m = reg_0_2&reg_0_4&reg_0_6&cdxi455m;
wire cdxi2089m = reg_0_2&reg_0_4&reg_0_5&cdxi394m;
wire cdxi2090m = reg_0_1&cdxi1501m;
wire cdxi2091m = reg_0_1&cdxi1502m;
wire cdxi2092m = reg_0_1&cdxi1503m;
wire cdxi2093m = reg_0_1&cdxi1504m;
wire cdxi2094m = reg_0_1&cdxi1505m;
wire cdxi2095m = reg_0_1&cdxi1506m;
wire cdxi2096m = reg_0_5&cdxi1006m;
wire cdxi2097m = reg_0_4&cdxi1043m;
wire cdxi2098m = reg_0_4&cdxi1044m;
wire cdxi2099m = reg_0_2&reg_0_6&cdxi456m;
wire cdxi2100m = reg_0_2&reg_0_5&cdxi475m;
wire cdxi2101m = reg_0_2&reg_0_4&cdxi1031m;
wire cdxi2102m = reg_0_1&cdxi1507m;
wire cdxi2103m = reg_0_1&cdxi1508m;
wire cdxi2104m = reg_0_1&cdxi1509m;
wire cdxi2105m = reg_0_1&cdxi1510m;
wire cdxi2106m = reg_0_6&cdxi1798m;
wire cdxi2107m = reg_0_5&cdxi995m;
wire cdxi2108m = reg_0_4&cdxi1032m;
wire cdxi2109m = reg_0_2&cdxi2079m;
wire cdxi2110m = reg_0_1&cdxi1496m;
wire cdxi2111m = (cdxi2081m ^ cdxi2082m ^ cdxi2083m ^ cdxi2084m ^ cdxi2085m ^ cdxi2086m ^ cdxi2087m ^ cdxi2088m ^ cdxi2089m ^ cdxi2090m ^ cdxi2091m ^ cdxi2092m ^ cdxi2093m ^ cdxi2094m ^ cdxi2095m ^ cdxi2096m ^ cdxi2097m ^ cdxi2098m ^ cdxi2099m ^ cdxi2100m ^ cdxi2101m ^ cdxi2102m ^ cdxi2103m ^ cdxi2104m ^ cdxi2105m ^ cdxi2106m ^ cdxi2107m ^ cdxi2108m ^ cdxi2109m ^ cdxi2110m ^ cdxi2080m);
wire cdxi2112m = reg_0_0&cdxi2111m;
wire cdxi2113m = cdxi363m&cdxi1268m ^ r106m;
wire cdxi2114m = cdxi977m&cdxi207m;
wire cdxi2115m = cdxi406m&cdxi657m;
wire cdxi2116m = cdxi363m&cdxi657m;
wire cdxi2117m = cdxi363m&cdxi562m;
wire cdxi2118m = cdxi977m&cdxi208m;
wire cdxi2119m = cdxi978m&cdxi271m;
wire cdxi2120m = cdxi363m&cdxi758m;
wire cdxi2121m = cdxi363m&cdxi759m;
wire cdxi2122m = cdxi363m&cdxi760m;
wire cdxi2123m = cdxi1268m&r7m;
wire cdxi2124m = cdxi1050m&r9m;
wire cdxi2125m = cdxi1339m&r11m;
wire cdxi2126m = cdxi977m&r12m;
wire cdxi2127m = cdxi385m&cdxi567m;
wire cdxi2128m = cdxi1124m&r16m;
wire cdxi2129m = cdxi978m&r17m;
wire cdxi2130m = cdxi363m&cdxi761m;
wire cdxi2131m = cdxi363m&cdxi762m;
wire cdxi2132m = cdxi363m&cdxi763m;
wire cdxi2133m = cdxi657m&r29m;
wire cdxi2134m = cdxi562m&r31m;
wire cdxi2135m = cdxi466m&r32m;
wire cdxi2136m = cdxi563m&r38m;
wire cdxi2137m = cdxi384m&r39m;
wire cdxi2138m = cdxi504m&r42m;
wire cdxi2139m = cdxi426m&r48m;
wire cdxi2140m = cdxi385m&r49m;
wire cdxi2141m = cdxi406m&r52m;
wire cdxi2142m = cdxi363m&r61m;
wire cdxi2143m = cdxi207m&r68m;
wire cdxi2144m = cdxi218m&r69m;
wire cdxi2145m = cdxi196m&r72m;
wire cdxi2146m = cdxi219m&r81m;
wire cdxi2147m = cdxi185m&r91m;
wire cdxi2148m = (cdxi2113m ^ cdxi2118m ^ cdxi2119m ^ cdxi2120m ^ cdxi2121m ^ cdxi2122m ^ cdxi2123m ^ cdxi2124m ^ cdxi2125m ^ cdxi2126m ^ cdxi2127m ^ cdxi2128m ^ cdxi2129m ^ cdxi2130m ^ cdxi2131m ^ cdxi2132m ^ cdxi2133m ^ cdxi2134m ^ cdxi2135m ^ cdxi2136m ^ cdxi2137m ^ cdxi2138m ^ cdxi2139m ^ cdxi2140m ^ cdxi2141m ^ cdxi2142m ^ cdxi2143m ^ cdxi2144m ^ cdxi2145m ^ cdxi2146m ^ cdxi2147m);
wire cdxi2149m = a0&cdxi2148m;
wire cdxi2150m = (reg_0_77);
wire cdxi2151m = (reg_0_99);
wire cdxi2152m = (reg_0_114);
wire cdxi2153m = reg_0_2&cdxi1286m;
wire cdxi2154m = reg_0_1&reg_0_4&reg_0_6&cdxi276m;
wire cdxi2155m = reg_0_1&reg_0_2&cdxi767m;
wire cdxi2156m = reg_0_1&reg_0_2&cdxi768m;
wire cdxi2157m = reg_0_1&reg_0_2&cdxi769m;
wire cdxi2158m = reg_0_4&cdxi1075m;
wire cdxi2159m = reg_0_2&cdxi1290m;
wire cdxi2160m = reg_0_2&cdxi1291m;
wire cdxi2161m = reg_0_2&cdxi1292m;
wire cdxi2162m = reg_0_1&reg_0_6&cdxi576m;
wire cdxi2163m = reg_0_1&reg_0_4&reg_0_7&cdxi224m;
wire cdxi2164m = reg_0_1&reg_0_4&reg_0_6&cdxi275m;
wire cdxi2165m = reg_0_1&reg_0_2&cdxi770m;
wire cdxi2166m = reg_0_1&reg_0_2&cdxi771m;
wire cdxi2167m = reg_0_1&reg_0_2&cdxi772m;
wire cdxi2168m = reg_0_6&reg_0_7&cdxi842m;
wire cdxi2169m = reg_0_4&cdxi1081m;
wire cdxi2170m = reg_0_4&cdxi1082m;
wire cdxi2171m = reg_0_2&cdxi1296m;
wire cdxi2172m = reg_0_2&cdxi1297m;
wire cdxi2173m = reg_0_2&cdxi1298m;
wire cdxi2174m = reg_0_1&reg_0_7&cdxi552m;
wire cdxi2175m = reg_0_1&reg_0_6&cdxi572m;
wire cdxi2176m = reg_0_1&reg_0_4&cdxi1069m;
wire cdxi2177m = reg_0_1&reg_0_2&cdxi766m;
wire cdxi2178m = reg_0_7&cdxi995m;
wire cdxi2179m = reg_0_6&cdxi2150m;
wire cdxi2180m = reg_0_4&cdxi1070m;
wire cdxi2181m = reg_0_2&cdxi1285m;
wire cdxi2182m = reg_0_1&cdxi2151m;
wire cdxi2183m = (cdxi2153m ^ cdxi2154m ^ cdxi2155m ^ cdxi2156m ^ cdxi2157m ^ cdxi2158m ^ cdxi2159m ^ cdxi2160m ^ cdxi2161m ^ cdxi2162m ^ cdxi2163m ^ cdxi2164m ^ cdxi2165m ^ cdxi2166m ^ cdxi2167m ^ cdxi2168m ^ cdxi2169m ^ cdxi2170m ^ cdxi2171m ^ cdxi2172m ^ cdxi2173m ^ cdxi2174m ^ cdxi2175m ^ cdxi2176m ^ cdxi2177m ^ cdxi2178m ^ cdxi2179m ^ cdxi2180m ^ cdxi2181m ^ cdxi2182m ^ cdxi2152m);
wire cdxi2184m = reg_0_0&cdxi2183m;
wire cdxi2185m = cdxi363m&cdxi1548m ^ r107m;
wire cdxi2186m = cdxi524m&cdxi657m;
wire cdxi2187m = cdxi446m&cdxi657m;
wire cdxi2188m = cdxi1013m&cdxi208m;
wire cdxi2189m = cdxi1014m&cdxi271m;
wire cdxi2190m = cdxi363m&cdxi658m;
wire cdxi2191m = cdxi363m&cdxi659m;
wire cdxi2192m = cdxi363m&cdxi660m;
wire cdxi2193m = cdxi1548m&r7m;
wire cdxi2194m = cdxi384m&cdxi489m;
wire cdxi2195m = cdxi1410m&r11m;
wire cdxi2196m = cdxi1013m&r12m;
wire cdxi2197m = cdxi385m&cdxi737m;
wire cdxi2198m = cdxi1161m&r16m;
wire cdxi2199m = cdxi1014m&r17m;
wire cdxi2200m = cdxi363m&cdxi661m;
wire cdxi2201m = cdxi363m&cdxi662m;
wire cdxi2202m = cdxi363m&cdxi663m;
wire cdxi2203m = cdxi657m&r30m;
wire cdxi2204m = cdxi485m&r31m;
wire cdxi2205m = cdxi638m&r32m;
wire cdxi2206m = cdxi563m&r40m;
wire cdxi2207m = cdxi384m&r41m;
wire cdxi2208m = cdxi524m&r42m;
wire cdxi2209m = cdxi426m&r50m;
wire cdxi2210m = cdxi385m&r51m;
wire cdxi2211m = cdxi446m&r52m;
wire cdxi2212m = cdxi363m&r62m;
wire cdxi2213m = cdxi207m&r70m;
wire cdxi2214m = cdxi218m&r71m;
wire cdxi2215m = cdxi240m&r72m;
wire cdxi2216m = cdxi219m&r82m;
wire cdxi2217m = cdxi185m&r92m;
wire cdxi2218m = (cdxi2185m ^ cdxi2188m ^ cdxi2189m ^ cdxi2190m ^ cdxi2191m ^ cdxi2192m ^ cdxi2193m ^ cdxi2194m ^ cdxi2195m ^ cdxi2196m ^ cdxi2197m ^ cdxi2198m ^ cdxi2199m ^ cdxi2200m ^ cdxi2201m ^ cdxi2202m ^ cdxi2203m ^ cdxi2204m ^ cdxi2205m ^ cdxi2206m ^ cdxi2207m ^ cdxi2208m ^ cdxi2209m ^ cdxi2210m ^ cdxi2211m ^ cdxi2212m ^ cdxi2213m ^ cdxi2214m ^ cdxi2215m ^ cdxi2216m ^ cdxi2217m);
wire cdxi2219m = a0&cdxi2218m;
wire cdxi2220m = (reg_0_90);
wire cdxi2221m = (reg_0_100);
wire cdxi2222m = (reg_0_115);
wire cdxi2223m = reg_0_2&reg_0_5&reg_0_6&cdxi213m;
wire cdxi2224m = reg_0_1&reg_0_5&reg_0_6&cdxi276m;
wire cdxi2225m = reg_0_1&reg_0_2&cdxi667m;
wire cdxi2226m = reg_0_1&reg_0_2&cdxi668m;
wire cdxi2227m = reg_0_1&reg_0_2&cdxi669m;
wire cdxi2228m = reg_0_5&cdxi1075m;
wire cdxi2229m = reg_0_2&reg_0_6&cdxi498m;
wire cdxi2230m = reg_0_2&reg_0_5&reg_0_7&cdxi394m;
wire cdxi2231m = reg_0_2&reg_0_5&reg_0_6&cdxi212m;
wire cdxi2232m = reg_0_1&reg_0_6&cdxi746m;
wire cdxi2233m = reg_0_1&reg_0_5&reg_0_7&cdxi224m;
wire cdxi2234m = reg_0_1&reg_0_5&reg_0_6&cdxi275m;
wire cdxi2235m = reg_0_1&reg_0_2&cdxi670m;
wire cdxi2236m = reg_0_1&reg_0_2&cdxi671m;
wire cdxi2237m = reg_0_1&reg_0_2&cdxi672m;
wire cdxi2238m = reg_0_6&reg_0_7&cdxi880m;
wire cdxi2239m = reg_0_5&cdxi1081m;
wire cdxi2240m = reg_0_5&cdxi1082m;
wire cdxi2241m = reg_0_2&reg_0_7&cdxi1031m;
wire cdxi2242m = reg_0_2&reg_0_6&cdxi494m;
wire cdxi2243m = reg_0_2&reg_0_5&cdxi1068m;
wire cdxi2244m = reg_0_1&reg_0_7&cdxi724m;
wire cdxi2245m = reg_0_1&reg_0_6&cdxi742m;
wire cdxi2246m = reg_0_1&reg_0_5&cdxi1069m;
wire cdxi2247m = reg_0_1&reg_0_2&cdxi666m;
wire cdxi2248m = reg_0_7&cdxi1032m;
wire cdxi2249m = reg_0_6&cdxi2010m;
wire cdxi2250m = reg_0_5&cdxi1070m;
wire cdxi2251m = reg_0_2&cdxi2220m;
wire cdxi2252m = reg_0_1&cdxi2221m;
wire cdxi2253m = (cdxi2223m ^ cdxi2224m ^ cdxi2225m ^ cdxi2226m ^ cdxi2227m ^ cdxi2228m ^ cdxi2229m ^ cdxi2230m ^ cdxi2231m ^ cdxi2232m ^ cdxi2233m ^ cdxi2234m ^ cdxi2235m ^ cdxi2236m ^ cdxi2237m ^ cdxi2238m ^ cdxi2239m ^ cdxi2240m ^ cdxi2241m ^ cdxi2242m ^ cdxi2243m ^ cdxi2244m ^ cdxi2245m ^ cdxi2246m ^ cdxi2247m ^ cdxi2248m ^ cdxi2249m ^ cdxi2250m ^ cdxi2251m ^ cdxi2252m ^ cdxi2222m);
wire cdxi2254m = reg_0_0&cdxi2253m;
wire cdxi2255m = cdxi362m&cdxi1479m ^ r108m;
wire cdxi2256m = cdxi405m&cdxi638m;
wire cdxi2257m = cdxi2256m&r0m;
wire cdxi2258m = cdxi1233m&cdxi291m;
wire cdxi2259m = cdxi362m&cdxi639m;
wire cdxi2260m = cdxi362m&cdxi640m;
wire cdxi2261m = cdxi362m&cdxi641m;
wire cdxi2262m = cdxi1479m&r8m;
wire cdxi2263m = cdxi582m&cdxi470m;
wire cdxi2264m = cdxi1088m&r10m;
wire cdxi2265m = cdxi1303m&r11m;
wire cdxi2266m = cdxi446m&cdxi605m;
wire cdxi2267m = cdxi978m&r19m;
wire cdxi2268m = cdxi1233m&r20m;
wire cdxi2269m = cdxi362m&cdxi642m;
wire cdxi2270m = cdxi362m&cdxi643m;
wire cdxi2271m = cdxi362m&cdxi644m;
wire cdxi2272m = cdxi638m&r33m;
wire cdxi2273m = cdxi466m&r34m;
wire cdxi2274m = cdxi445m&r35m;
wire cdxi2275m = cdxi601m&r37m;
wire cdxi2276m = cdxi582m&r38m;
wire cdxi2277m = cdxi405m&r40m;
wire cdxi2278m = cdxi385m&r53m;
wire cdxi2279m = cdxi446m&r54m;
wire cdxi2280m = cdxi406m&r56m;
wire cdxi2281m = cdxi362m&r59m;
wire cdxi2282m = cdxi218m&r73m;
wire cdxi2283m = cdxi240m&r74m;
wire cdxi2284m = cdxi196m&r76m;
wire cdxi2285m = cdxi184m&r79m;
wire cdxi2286m = cdxi185m&r93m;
wire cdxi2287m = (cdxi2255m ^ cdxi2257m ^ cdxi2258m ^ cdxi2259m ^ cdxi2260m ^ cdxi2261m ^ cdxi2262m ^ cdxi2263m ^ cdxi2264m ^ cdxi2265m ^ cdxi2266m ^ cdxi2267m ^ cdxi2268m ^ cdxi2269m ^ cdxi2270m ^ cdxi2271m ^ cdxi2272m ^ cdxi2273m ^ cdxi2274m ^ cdxi2275m ^ cdxi2276m ^ cdxi2277m ^ cdxi2278m ^ cdxi2279m ^ cdxi2280m ^ cdxi2281m ^ cdxi2282m ^ cdxi2283m ^ cdxi2284m ^ cdxi2285m ^ cdxi2286m);
wire cdxi2288m = a0&cdxi2287m;
wire cdxi2289m = (reg_0_116);
wire cdxi2290m = reg_0_3&reg_0_4&reg_0_5&reg_0_6&cdxi130m;
wire cdxi2291m = reg_0_1&cdxi1704m;
wire cdxi2292m = reg_0_1&cdxi1705m;
wire cdxi2293m = reg_0_1&cdxi1706m;
wire cdxi2294m = reg_0_1&cdxi1707m;
wire cdxi2295m = reg_0_4&reg_0_5&reg_0_6&cdxi190m;
wire cdxi2296m = reg_0_3&reg_0_5&cdxi479m;
wire cdxi2297m = reg_0_3&reg_0_4&reg_0_6&cdxi455m;
wire cdxi2298m = reg_0_3&reg_0_4&reg_0_5&cdxi394m;
wire cdxi2299m = reg_0_1&cdxi1708m;
wire cdxi2300m = reg_0_1&cdxi1709m;
wire cdxi2301m = reg_0_1&cdxi1710m;
wire cdxi2302m = reg_0_1&cdxi1711m;
wire cdxi2303m = reg_0_1&cdxi1712m;
wire cdxi2304m = reg_0_1&cdxi1713m;
wire cdxi2305m = reg_0_5&cdxi1116m;
wire cdxi2306m = reg_0_4&reg_0_6&cdxi881m;
wire cdxi2307m = reg_0_4&reg_0_5&cdxi919m;
wire cdxi2308m = reg_0_3&reg_0_6&cdxi456m;
wire cdxi2309m = reg_0_3&reg_0_5&cdxi475m;
wire cdxi2310m = reg_0_3&reg_0_4&cdxi1031m;
wire cdxi2311m = reg_0_1&cdxi1714m;
wire cdxi2312m = reg_0_1&cdxi1715m;
wire cdxi2313m = reg_0_1&cdxi1716m;
wire cdxi2314m = reg_0_1&cdxi1717m;
wire cdxi2315m = reg_0_6&cdxi1799m;
wire cdxi2316m = reg_0_5&cdxi1105m;
wire cdxi2317m = reg_0_4&cdxi1939m;
wire cdxi2318m = reg_0_3&cdxi2079m;
wire cdxi2319m = reg_0_1&cdxi1703m;
wire cdxi2320m = (cdxi2290m ^ cdxi2291m ^ cdxi2292m ^ cdxi2293m ^ cdxi2294m ^ cdxi2295m ^ cdxi2296m ^ cdxi2297m ^ cdxi2298m ^ cdxi2299m ^ cdxi2300m ^ cdxi2301m ^ cdxi2302m ^ cdxi2303m ^ cdxi2304m ^ cdxi2305m ^ cdxi2306m ^ cdxi2307m ^ cdxi2308m ^ cdxi2309m ^ cdxi2310m ^ cdxi2311m ^ cdxi2312m ^ cdxi2313m ^ cdxi2314m ^ cdxi2315m ^ cdxi2316m ^ cdxi2317m ^ cdxi2318m ^ cdxi2319m ^ cdxi2289m);
wire cdxi2321m = reg_0_0&cdxi2320m;
wire cdxi2322m = cdxi362m&cdxi1232m ^ r109m;
wire cdxi2323m = cdxi405m&cdxi485m;
wire cdxi2324m = cdxi406m&cdxi485m;
wire cdxi2325m = cdxi362m&cdxi562m;
wire cdxi2326m = cdxi405m&cdxi486m;
wire cdxi2327m = cdxi406m&cdxi620m;
wire cdxi2328m = cdxi362m&cdxi802m;
wire cdxi2329m = cdxi362m&cdxi803m;
wire cdxi2330m = cdxi362m&cdxi804m;
wire cdxi2331m = cdxi445m&cdxi430m;
wire cdxi2332m = cdxi1160m&r9m;
wire cdxi2333m = cdxi405m&cdxi489m;
wire cdxi2334m = cdxi405m&cdxi490m;
wire cdxi2335m = cdxi446m&cdxi781m;
wire cdxi2336m = cdxi406m&cdxi623m;
wire cdxi2337m = cdxi406m&cdxi624m;
wire cdxi2338m = cdxi362m&cdxi805m;
wire cdxi2339m = cdxi362m&cdxi806m;
wire cdxi2340m = cdxi362m&cdxi807m;
wire cdxi2341m = cdxi485m&r33m;
wire cdxi2342m = cdxi562m&r34m;
wire cdxi2343m = cdxi445m&r36m;
wire cdxi2344m = cdxi425m&r37m;
wire cdxi2345m = cdxi582m&r39m;
wire cdxi2346m = cdxi405m&r41m;
wire cdxi2347m = cdxi426m&r53m;
wire cdxi2348m = cdxi446m&r55m;
wire cdxi2349m = cdxi406m&r57m;
wire cdxi2350m = cdxi362m&r60m;
wire cdxi2351m = cdxi207m&r73m;
wire cdxi2352m = cdxi240m&r75m;
wire cdxi2353m = cdxi196m&r77m;
wire cdxi2354m = cdxi184m&r80m;
wire cdxi2355m = cdxi185m&r94m;
wire cdxi2356m = (cdxi2322m ^ cdxi2326m ^ cdxi2327m ^ cdxi2328m ^ cdxi2329m ^ cdxi2330m ^ cdxi2331m ^ cdxi2332m ^ cdxi2333m ^ cdxi2334m ^ cdxi2335m ^ cdxi2336m ^ cdxi2337m ^ cdxi2338m ^ cdxi2339m ^ cdxi2340m ^ cdxi2341m ^ cdxi2342m ^ cdxi2343m ^ cdxi2344m ^ cdxi2345m ^ cdxi2346m ^ cdxi2347m ^ cdxi2348m ^ cdxi2349m ^ cdxi2350m ^ cdxi2351m ^ cdxi2352m ^ cdxi2353m ^ cdxi2354m ^ cdxi2355m);
wire cdxi2357m = a0&cdxi2356m;
wire cdxi2358m = (reg_0_117);
wire cdxi2359m = reg_0_3&cdxi1251m;
wire cdxi2360m = reg_0_1&cdxi1636m;
wire cdxi2361m = reg_0_1&cdxi1637m;
wire cdxi2362m = reg_0_1&cdxi1638m;
wire cdxi2363m = reg_0_1&cdxi1639m;
wire cdxi2364m = reg_0_4&cdxi1183m;
wire cdxi2365m = reg_0_3&cdxi1255m;
wire cdxi2366m = reg_0_3&cdxi1256m;
wire cdxi2367m = reg_0_3&cdxi1257m;
wire cdxi2368m = reg_0_1&cdxi1640m;
wire cdxi2369m = reg_0_1&cdxi1641m;
wire cdxi2370m = reg_0_1&cdxi1642m;
wire cdxi2371m = reg_0_1&cdxi1643m;
wire cdxi2372m = reg_0_1&cdxi1644m;
wire cdxi2373m = reg_0_1&cdxi1645m;
wire cdxi2374m = reg_0_5&cdxi1153m;
wire cdxi2375m = reg_0_4&cdxi1189m;
wire cdxi2376m = reg_0_4&cdxi1190m;
wire cdxi2377m = reg_0_3&cdxi1261m;
wire cdxi2378m = reg_0_3&cdxi1262m;
wire cdxi2379m = reg_0_3&cdxi1263m;
wire cdxi2380m = reg_0_1&cdxi1646m;
wire cdxi2381m = reg_0_1&cdxi1647m;
wire cdxi2382m = reg_0_1&cdxi1648m;
wire cdxi2383m = reg_0_1&cdxi1649m;
wire cdxi2384m = reg_0_7&cdxi1799m;
wire cdxi2385m = reg_0_5&cdxi1142m;
wire cdxi2386m = reg_0_4&cdxi1178m;
wire cdxi2387m = reg_0_3&cdxi1250m;
wire cdxi2388m = reg_0_1&cdxi1635m;
wire cdxi2389m = (cdxi2359m ^ cdxi2360m ^ cdxi2361m ^ cdxi2362m ^ cdxi2363m ^ cdxi2364m ^ cdxi2365m ^ cdxi2366m ^ cdxi2367m ^ cdxi2368m ^ cdxi2369m ^ cdxi2370m ^ cdxi2371m ^ cdxi2372m ^ cdxi2373m ^ cdxi2374m ^ cdxi2375m ^ cdxi2376m ^ cdxi2377m ^ cdxi2378m ^ cdxi2379m ^ cdxi2380m ^ cdxi2381m ^ cdxi2382m ^ cdxi2383m ^ cdxi2384m ^ cdxi2385m ^ cdxi2386m ^ cdxi2387m ^ cdxi2388m ^ cdxi2358m);
wire cdxi2390m = reg_0_0&cdxi2389m;
wire cdxi2391m = cdxi406m&cdxi1548m ^ r112m;
wire cdxi2392m = cdxi445m&cdxi657m;
wire cdxi2393m = cdxi1479m&cdxi208m;
wire cdxi2394m = cdxi446m&cdxi758m;
wire cdxi2395m = cdxi406m&cdxi658m;
wire cdxi2396m = cdxi406m&cdxi659m;
wire cdxi2397m = cdxi406m&cdxi660m;
wire cdxi2398m = cdxi1548m&r9m;
wire cdxi2399m = cdxi466m&cdxi489m;
wire cdxi2400m = cdxi1232m&r11m;
wire cdxi2401m = cdxi1479m&r12m;
wire cdxi2402m = cdxi385m&cdxi805m;
wire cdxi2403m = cdxi446m&cdxi761m;
wire cdxi2404m = cdxi446m&cdxi762m;
wire cdxi2405m = cdxi406m&cdxi661m;
wire cdxi2406m = cdxi406m&cdxi662m;
wire cdxi2407m = cdxi406m&cdxi663m;
wire cdxi2408m = cdxi657m&r37m;
wire cdxi2409m = cdxi485m&r38m;
wire cdxi2410m = cdxi638m&r39m;
wire cdxi2411m = cdxi562m&r40m;
wire cdxi2412m = cdxi466m&r41m;
wire cdxi2413m = cdxi445m&r42m;
wire cdxi2414m = cdxi426m&r59m;
wire cdxi2415m = cdxi385m&r60m;
wire cdxi2416m = cdxi446m&r61m;
wire cdxi2417m = cdxi406m&r62m;
wire cdxi2418m = cdxi207m&r79m;
wire cdxi2419m = cdxi218m&r80m;
wire cdxi2420m = cdxi240m&r81m;
wire cdxi2421m = cdxi196m&r82m;
wire cdxi2422m = cdxi185m&r97m;
wire cdxi2423m = (cdxi2391m ^ cdxi2393m ^ cdxi2394m ^ cdxi2395m ^ cdxi2396m ^ cdxi2397m ^ cdxi2398m ^ cdxi2399m ^ cdxi2400m ^ cdxi2401m ^ cdxi2402m ^ cdxi2403m ^ cdxi2404m ^ cdxi2405m ^ cdxi2406m ^ cdxi2407m ^ cdxi2408m ^ cdxi2409m ^ cdxi2410m ^ cdxi2411m ^ cdxi2412m ^ cdxi2413m ^ cdxi2414m ^ cdxi2415m ^ cdxi2416m ^ cdxi2417m ^ cdxi2418m ^ cdxi2419m ^ cdxi2420m ^ cdxi2421m ^ cdxi2422m);
wire cdxi2424m = a0&cdxi2423m;
wire cdxi2425m = (reg_0_120);
wire cdxi2426m = reg_0_4&reg_0_5&reg_0_6&cdxi213m;
wire cdxi2427m = reg_0_1&cdxi1744m;
wire cdxi2428m = reg_0_1&cdxi1745m;
wire cdxi2429m = reg_0_1&cdxi1746m;
wire cdxi2430m = reg_0_1&cdxi1747m;
wire cdxi2431m = reg_0_5&cdxi1290m;
wire cdxi2432m = reg_0_4&reg_0_6&cdxi498m;
wire cdxi2433m = reg_0_4&reg_0_5&reg_0_7&cdxi394m;
wire cdxi2434m = reg_0_4&reg_0_5&reg_0_6&cdxi212m;
wire cdxi2435m = reg_0_1&cdxi1748m;
wire cdxi2436m = reg_0_1&cdxi1749m;
wire cdxi2437m = reg_0_1&cdxi1750m;
wire cdxi2438m = reg_0_1&cdxi1751m;
wire cdxi2439m = reg_0_1&cdxi1752m;
wire cdxi2440m = reg_0_1&cdxi1753m;
wire cdxi2441m = reg_0_6&cdxi1261m;
wire cdxi2442m = reg_0_5&cdxi1296m;
wire cdxi2443m = reg_0_5&cdxi1297m;
wire cdxi2444m = reg_0_4&reg_0_7&cdxi1031m;
wire cdxi2445m = reg_0_4&reg_0_6&cdxi494m;
wire cdxi2446m = reg_0_4&reg_0_5&cdxi1068m;
wire cdxi2447m = reg_0_1&cdxi1754m;
wire cdxi2448m = reg_0_1&cdxi1755m;
wire cdxi2449m = reg_0_1&cdxi1756m;
wire cdxi2450m = reg_0_1&cdxi1757m;
wire cdxi2451m = reg_0_7&cdxi2079m;
wire cdxi2452m = reg_0_6&cdxi1250m;
wire cdxi2453m = reg_0_5&cdxi1285m;
wire cdxi2454m = reg_0_4&cdxi2220m;
wire cdxi2455m = reg_0_1&cdxi1743m;
wire cdxi2456m = (cdxi2426m ^ cdxi2427m ^ cdxi2428m ^ cdxi2429m ^ cdxi2430m ^ cdxi2431m ^ cdxi2432m ^ cdxi2433m ^ cdxi2434m ^ cdxi2435m ^ cdxi2436m ^ cdxi2437m ^ cdxi2438m ^ cdxi2439m ^ cdxi2440m ^ cdxi2441m ^ cdxi2442m ^ cdxi2443m ^ cdxi2444m ^ cdxi2445m ^ cdxi2446m ^ cdxi2447m ^ cdxi2448m ^ cdxi2449m ^ cdxi2450m ^ cdxi2451m ^ cdxi2452m ^ cdxi2453m ^ cdxi2454m ^ cdxi2455m ^ cdxi2425m);
wire cdxi2457m = reg_0_0&cdxi2456m;
wire cdxi2458m = cdxi361m&cdxi1232m ^ r114m;
wire cdxi2459m = cdxi219m&cdxi1232m;
wire cdxi2460m = cdxi361m&cdxi562m;
wire cdxi2461m = cdxi405m&cdxi734m;
wire cdxi2462m = cdxi1304m&cdxi230m;
wire cdxi2463m = cdxi361m&cdxi802m;
wire cdxi2464m = cdxi361m&cdxi803m;
wire cdxi2465m = cdxi361m&cdxi804m;
wire cdxi2466m = cdxi1232m&r13m;
wire cdxi2467m = cdxi1160m&r14m;
wire cdxi2468m = cdxi405m&cdxi737m;
wire cdxi2469m = cdxi405m&cdxi738m;
wire cdxi2470m = cdxi1410m&r18m;
wire cdxi2471m = cdxi504m&cdxi623m;
wire cdxi2472m = cdxi1304m&r21m;
wire cdxi2473m = cdxi361m&cdxi805m;
wire cdxi2474m = cdxi361m&cdxi806m;
wire cdxi2475m = cdxi361m&cdxi807m;
wire cdxi2476m = cdxi485m&r43m;
wire cdxi2477m = cdxi562m&r44m;
wire cdxi2478m = cdxi445m&r46m;
wire cdxi2479m = cdxi425m&r47m;
wire cdxi2480m = cdxi582m&r49m;
wire cdxi2481m = cdxi405m&r51m;
wire cdxi2482m = cdxi563m&r53m;
wire cdxi2483m = cdxi524m&r55m;
wire cdxi2484m = cdxi504m&r57m;
wire cdxi2485m = cdxi361m&r60m;
wire cdxi2486m = cdxi207m&r83m;
wire cdxi2487m = cdxi240m&r85m;
wire cdxi2488m = cdxi196m&r87m;
wire cdxi2489m = cdxi184m&r90m;
wire cdxi2490m = cdxi219m&r94m;
wire cdxi2491m = (cdxi2458m ^ cdxi2461m ^ cdxi2462m ^ cdxi2463m ^ cdxi2464m ^ cdxi2465m ^ cdxi2466m ^ cdxi2467m ^ cdxi2468m ^ cdxi2469m ^ cdxi2470m ^ cdxi2471m ^ cdxi2472m ^ cdxi2473m ^ cdxi2474m ^ cdxi2475m ^ cdxi2476m ^ cdxi2477m ^ cdxi2478m ^ cdxi2479m ^ cdxi2480m ^ cdxi2481m ^ cdxi2482m ^ cdxi2483m ^ cdxi2484m ^ cdxi2485m ^ cdxi2486m ^ cdxi2487m ^ cdxi2488m ^ cdxi2489m ^ cdxi2490m);
wire cdxi2492m = a0&cdxi2491m;
wire cdxi2493m = (reg_0_122);
wire cdxi2494m = reg_0_3&cdxi1531m;
wire cdxi2495m = reg_0_2&cdxi1636m;
wire cdxi2496m = reg_0_2&cdxi1637m;
wire cdxi2497m = reg_0_2&cdxi1638m;
wire cdxi2498m = reg_0_2&cdxi1639m;
wire cdxi2499m = reg_0_4&cdxi1432m;
wire cdxi2500m = reg_0_3&cdxi1535m;
wire cdxi2501m = reg_0_3&cdxi1536m;
wire cdxi2502m = reg_0_3&cdxi1537m;
wire cdxi2503m = reg_0_2&cdxi1640m;
wire cdxi2504m = reg_0_2&cdxi1641m;
wire cdxi2505m = reg_0_2&cdxi1642m;
wire cdxi2506m = reg_0_2&cdxi1643m;
wire cdxi2507m = reg_0_2&cdxi1644m;
wire cdxi2508m = reg_0_2&cdxi1645m;
wire cdxi2509m = reg_0_5&cdxi1367m;
wire cdxi2510m = reg_0_4&cdxi1438m;
wire cdxi2511m = reg_0_4&cdxi1439m;
wire cdxi2512m = reg_0_3&cdxi1541m;
wire cdxi2513m = reg_0_3&cdxi1542m;
wire cdxi2514m = reg_0_3&cdxi1543m;
wire cdxi2515m = reg_0_2&cdxi1646m;
wire cdxi2516m = reg_0_2&cdxi1647m;
wire cdxi2517m = reg_0_2&cdxi1648m;
wire cdxi2518m = reg_0_2&cdxi1649m;
wire cdxi2519m = reg_0_7&cdxi1321m;
wire cdxi2520m = reg_0_5&cdxi1356m;
wire cdxi2521m = reg_0_4&cdxi1427m;
wire cdxi2522m = reg_0_3&cdxi1530m;
wire cdxi2523m = reg_0_2&cdxi1635m;
wire cdxi2524m = (cdxi2494m ^ cdxi2495m ^ cdxi2496m ^ cdxi2497m ^ cdxi2498m ^ cdxi2499m ^ cdxi2500m ^ cdxi2501m ^ cdxi2502m ^ cdxi2503m ^ cdxi2504m ^ cdxi2505m ^ cdxi2506m ^ cdxi2507m ^ cdxi2508m ^ cdxi2509m ^ cdxi2510m ^ cdxi2511m ^ cdxi2512m ^ cdxi2513m ^ cdxi2514m ^ cdxi2515m ^ cdxi2516m ^ cdxi2517m ^ cdxi2518m ^ cdxi2519m ^ cdxi2520m ^ cdxi2521m ^ cdxi2522m ^ cdxi2523m ^ cdxi2493m);
wire cdxi2525m = reg_0_0&cdxi2524m;
wire cdxi2526m = cdxi361m&cdxi1268m ^ r115m;
wire cdxi2527m = cdxi405m&cdxi657m;
wire cdxi2528m = cdxi361m&cdxi657m;
wire cdxi2529m = cdxi1088m&cdxi271m;
wire cdxi2530m = cdxi977m&cdxi230m;
wire cdxi2531m = cdxi361m&cdxi758m;
wire cdxi2532m = cdxi361m&cdxi759m;
wire cdxi2533m = cdxi361m&cdxi760m;
wire cdxi2534m = cdxi1268m&r13m;
wire cdxi2535m = cdxi601m&cdxi567m;
wire cdxi2536m = cdxi1123m&r16m;
wire cdxi2537m = cdxi1088m&r17m;
wire cdxi2538m = cdxi384m&cdxi781m;
wire cdxi2539m = cdxi1339m&r20m;
wire cdxi2540m = cdxi977m&r21m;
wire cdxi2541m = cdxi361m&cdxi761m;
wire cdxi2542m = cdxi361m&cdxi762m;
wire cdxi2543m = cdxi361m&cdxi763m;
wire cdxi2544m = cdxi657m&r43m;
wire cdxi2545m = cdxi562m&r45m;
wire cdxi2546m = cdxi466m&r46m;
wire cdxi2547m = cdxi425m&r48m;
wire cdxi2548m = cdxi601m&r49m;
wire cdxi2549m = cdxi405m&r52m;
wire cdxi2550m = cdxi563m&r54m;
wire cdxi2551m = cdxi384m&r55m;
wire cdxi2552m = cdxi504m&r58m;
wire cdxi2553m = cdxi361m&r61m;
wire cdxi2554m = cdxi207m&r84m;
wire cdxi2555m = cdxi218m&r85m;
wire cdxi2556m = cdxi196m&r88m;
wire cdxi2557m = cdxi184m&r91m;
wire cdxi2558m = cdxi219m&r95m;
wire cdxi2559m = (cdxi2526m ^ cdxi2529m ^ cdxi2530m ^ cdxi2531m ^ cdxi2532m ^ cdxi2533m ^ cdxi2534m ^ cdxi2535m ^ cdxi2536m ^ cdxi2537m ^ cdxi2538m ^ cdxi2539m ^ cdxi2540m ^ cdxi2541m ^ cdxi2542m ^ cdxi2543m ^ cdxi2544m ^ cdxi2545m ^ cdxi2546m ^ cdxi2547m ^ cdxi2548m ^ cdxi2549m ^ cdxi2550m ^ cdxi2551m ^ cdxi2552m ^ cdxi2553m ^ cdxi2554m ^ cdxi2555m ^ cdxi2556m ^ cdxi2557m ^ cdxi2558m);
wire cdxi2560m = a0&cdxi2559m;
wire cdxi2561m = (reg_0_123);
wire cdxi2562m = reg_0_3&reg_0_4&reg_0_6&cdxi276m;
wire cdxi2563m = reg_0_2&cdxi1670m;
wire cdxi2564m = reg_0_2&cdxi1671m;
wire cdxi2565m = reg_0_2&cdxi1672m;
wire cdxi2566m = reg_0_2&cdxi1673m;
wire cdxi2567m = reg_0_4&cdxi1466m;
wire cdxi2568m = reg_0_3&reg_0_6&cdxi576m;
wire cdxi2569m = reg_0_3&reg_0_4&reg_0_7&cdxi224m;
wire cdxi2570m = reg_0_3&reg_0_4&reg_0_6&cdxi275m;
wire cdxi2571m = reg_0_2&cdxi1674m;
wire cdxi2572m = reg_0_2&cdxi1675m;
wire cdxi2573m = reg_0_2&cdxi1676m;
wire cdxi2574m = reg_0_2&cdxi1677m;
wire cdxi2575m = reg_0_2&cdxi1678m;
wire cdxi2576m = reg_0_2&cdxi1679m;
wire cdxi2577m = reg_0_6&cdxi1367m;
wire cdxi2578m = reg_0_4&cdxi1472m;
wire cdxi2579m = reg_0_4&cdxi1473m;
wire cdxi2580m = reg_0_3&reg_0_7&cdxi552m;
wire cdxi2581m = reg_0_3&reg_0_6&cdxi572m;
wire cdxi2582m = reg_0_3&reg_0_4&cdxi1069m;
wire cdxi2583m = reg_0_2&cdxi1680m;
wire cdxi2584m = reg_0_2&cdxi1681m;
wire cdxi2585m = reg_0_2&cdxi1682m;
wire cdxi2586m = reg_0_2&cdxi1683m;
wire cdxi2587m = reg_0_7&cdxi1599m;
wire cdxi2588m = reg_0_6&cdxi1356m;
wire cdxi2589m = reg_0_4&cdxi1461m;
wire cdxi2590m = reg_0_3&cdxi2151m;
wire cdxi2591m = reg_0_2&cdxi1669m;
wire cdxi2592m = (cdxi2562m ^ cdxi2563m ^ cdxi2564m ^ cdxi2565m ^ cdxi2566m ^ cdxi2567m ^ cdxi2568m ^ cdxi2569m ^ cdxi2570m ^ cdxi2571m ^ cdxi2572m ^ cdxi2573m ^ cdxi2574m ^ cdxi2575m ^ cdxi2576m ^ cdxi2577m ^ cdxi2578m ^ cdxi2579m ^ cdxi2580m ^ cdxi2581m ^ cdxi2582m ^ cdxi2583m ^ cdxi2584m ^ cdxi2585m ^ cdxi2586m ^ cdxi2587m ^ cdxi2588m ^ cdxi2589m ^ cdxi2590m ^ cdxi2591m ^ cdxi2561m);
wire cdxi2593m = reg_0_0&cdxi2592m;
wire cdxi2594m = cdxi1304m&cdxi657m ^ r117m;
wire cdxi2595m = cdxi1479m&cdxi271m;
wire cdxi2596m = cdxi524m&cdxi758m;
wire cdxi2597m = cdxi977m&cdxi261m;
wire cdxi2598m = cdxi1304m&cdxi337m;
wire cdxi2599m = cdxi1304m&cdxi338m;
wire cdxi2600m = cdxi638m&cdxi567m;
wire cdxi2601m = cdxi466m&cdxi737m;
wire cdxi2602m = cdxi1232m&r16m;
wire cdxi2603m = cdxi1479m&r17m;
wire cdxi2604m = cdxi384m&cdxi805m;
wire cdxi2605m = cdxi1410m&r23m;
wire cdxi2606m = cdxi524m&cdxi762m;
wire cdxi2607m = cdxi504m&cdxi661m;
wire cdxi2608m = cdxi977m&r26m;
wire cdxi2609m = cdxi1304m&r27m;
wire cdxi2610m = cdxi657m&r47m;
wire cdxi2611m = cdxi485m&r48m;
wire cdxi2612m = cdxi638m&r49m;
wire cdxi2613m = cdxi562m&r50m;
wire cdxi2614m = cdxi466m&r51m;
wire cdxi2615m = cdxi445m&r52m;
wire cdxi2616m = cdxi563m&r59m;
wire cdxi2617m = cdxi384m&r60m;
wire cdxi2618m = cdxi524m&r61m;
wire cdxi2619m = cdxi504m&r62m;
wire cdxi2620m = cdxi207m&r89m;
wire cdxi2621m = cdxi218m&r90m;
wire cdxi2622m = cdxi240m&r91m;
wire cdxi2623m = cdxi196m&r92m;
wire cdxi2624m = cdxi219m&r97m;
wire cdxi2625m = (cdxi2594m ^ cdxi2595m ^ cdxi2596m ^ cdxi2597m ^ cdxi2598m ^ cdxi2599m ^ cdxi2600m ^ cdxi2601m ^ cdxi2602m ^ cdxi2603m ^ cdxi2604m ^ cdxi2605m ^ cdxi2606m ^ cdxi2607m ^ cdxi2608m ^ cdxi2609m ^ cdxi2610m ^ cdxi2611m ^ cdxi2612m ^ cdxi2613m ^ cdxi2614m ^ cdxi2615m ^ cdxi2616m ^ cdxi2617m ^ cdxi2618m ^ cdxi2619m ^ cdxi2620m ^ cdxi2621m ^ cdxi2622m ^ cdxi2623m ^ cdxi2624m);
wire cdxi2626m = a0&cdxi2625m;
wire cdxi2627m = (reg_0_125);
wire cdxi2628m = reg_0_4&reg_0_5&reg_0_6&cdxi276m;
wire cdxi2629m = reg_0_2&cdxi1744m;
wire cdxi2630m = reg_0_2&cdxi1745m;
wire cdxi2631m = reg_0_2&cdxi1746m;
wire cdxi2632m = reg_0_2&cdxi1747m;
wire cdxi2633m = reg_0_5&reg_0_6&cdxi576m;
wire cdxi2634m = reg_0_4&reg_0_6&cdxi746m;
wire cdxi2635m = reg_0_4&reg_0_5&reg_0_7&cdxi224m;
wire cdxi2636m = reg_0_4&reg_0_5&reg_0_6&cdxi275m;
wire cdxi2637m = reg_0_2&cdxi1748m;
wire cdxi2638m = reg_0_2&cdxi1749m;
wire cdxi2639m = reg_0_2&cdxi1750m;
wire cdxi2640m = reg_0_2&cdxi1751m;
wire cdxi2641m = reg_0_2&cdxi1752m;
wire cdxi2642m = reg_0_2&cdxi1753m;
wire cdxi2643m = reg_0_6&cdxi1541m;
wire cdxi2644m = reg_0_5&reg_0_7&cdxi552m;
wire cdxi2645m = reg_0_5&reg_0_6&cdxi572m;
wire cdxi2646m = reg_0_4&reg_0_7&cdxi724m;
wire cdxi2647m = reg_0_4&reg_0_6&cdxi742m;
wire cdxi2648m = reg_0_4&reg_0_5&cdxi1069m;
wire cdxi2649m = reg_0_2&cdxi1754m;
wire cdxi2650m = reg_0_2&cdxi1755m;
wire cdxi2651m = reg_0_2&cdxi1756m;
wire cdxi2652m = reg_0_2&cdxi1757m;
wire cdxi2653m = reg_0_7&cdxi1496m;
wire cdxi2654m = reg_0_6&cdxi1530m;
wire cdxi2655m = reg_0_5&cdxi2151m;
wire cdxi2656m = reg_0_4&cdxi2221m;
wire cdxi2657m = reg_0_2&cdxi1743m;
wire cdxi2658m = (cdxi2628m ^ cdxi2629m ^ cdxi2630m ^ cdxi2631m ^ cdxi2632m ^ cdxi2633m ^ cdxi2634m ^ cdxi2635m ^ cdxi2636m ^ cdxi2637m ^ cdxi2638m ^ cdxi2639m ^ cdxi2640m ^ cdxi2641m ^ cdxi2642m ^ cdxi2643m ^ cdxi2644m ^ cdxi2645m ^ cdxi2646m ^ cdxi2647m ^ cdxi2648m ^ cdxi2649m ^ cdxi2650m ^ cdxi2651m ^ cdxi2652m ^ cdxi2653m ^ cdxi2654m ^ cdxi2655m ^ cdxi2656m ^ cdxi2657m ^ cdxi2627m);
wire cdxi2659m = reg_0_0&cdxi2658m;
wire cdxi2660m = cdxi405m&cdxi1548m ^ r118m;
wire cdxi2661m = cdxi582m&cdxi657m;
wire cdxi2662m = cdxi1479m&cdxi230m;
wire cdxi2663m = cdxi582m&cdxi758m;
wire cdxi2664m = cdxi405m&cdxi658m;
wire cdxi2665m = cdxi405m&cdxi659m;
wire cdxi2666m = cdxi405m&cdxi660m;
wire cdxi2667m = cdxi638m&cdxi781m;
wire cdxi2668m = cdxi466m&cdxi623m;
wire cdxi2669m = cdxi1232m&r20m;
wire cdxi2670m = cdxi1479m&r21m;
wire cdxi2671m = cdxi601m&cdxi805m;
wire cdxi2672m = cdxi1160m&r23m;
wire cdxi2673m = cdxi582m&cdxi762m;
wire cdxi2674m = cdxi405m&cdxi661m;
wire cdxi2675m = cdxi405m&cdxi662m;
wire cdxi2676m = cdxi405m&cdxi663m;
wire cdxi2677m = cdxi657m&r53m;
wire cdxi2678m = cdxi485m&r54m;
wire cdxi2679m = cdxi638m&r55m;
wire cdxi2680m = cdxi562m&r56m;
wire cdxi2681m = cdxi466m&r57m;
wire cdxi2682m = cdxi445m&r58m;
wire cdxi2683m = cdxi425m&r59m;
wire cdxi2684m = cdxi601m&r60m;
wire cdxi2685m = cdxi582m&r61m;
wire cdxi2686m = cdxi405m&r62m;
wire cdxi2687m = cdxi207m&r93m;
wire cdxi2688m = cdxi218m&r94m;
wire cdxi2689m = cdxi240m&r95m;
wire cdxi2690m = cdxi196m&r96m;
wire cdxi2691m = cdxi184m&r97m;
wire cdxi2692m = (cdxi2660m ^ cdxi2662m ^ cdxi2663m ^ cdxi2664m ^ cdxi2665m ^ cdxi2666m ^ cdxi2667m ^ cdxi2668m ^ cdxi2669m ^ cdxi2670m ^ cdxi2671m ^ cdxi2672m ^ cdxi2673m ^ cdxi2674m ^ cdxi2675m ^ cdxi2676m ^ cdxi2677m ^ cdxi2678m ^ cdxi2679m ^ cdxi2680m ^ cdxi2681m ^ cdxi2682m ^ cdxi2683m ^ cdxi2684m ^ cdxi2685m ^ cdxi2686m ^ cdxi2687m ^ cdxi2688m ^ cdxi2689m ^ cdxi2690m ^ cdxi2691m);
wire cdxi2693m = a0&cdxi2692m;
wire cdxi2694m = (reg_0_126);
wire cdxi2695m = reg_0_4&cdxi1566m;
wire cdxi2696m = reg_0_3&cdxi1744m;
wire cdxi2697m = reg_0_3&cdxi1745m;
wire cdxi2698m = reg_0_3&cdxi1746m;
wire cdxi2699m = reg_0_3&cdxi1747m;
wire cdxi2700m = reg_0_5&cdxi1674m;
wire cdxi2701m = reg_0_4&cdxi1570m;
wire cdxi2702m = reg_0_4&cdxi1571m;
wire cdxi2703m = reg_0_4&cdxi1572m;
wire cdxi2704m = reg_0_3&cdxi1748m;
wire cdxi2705m = reg_0_3&cdxi1749m;
wire cdxi2706m = reg_0_3&cdxi1750m;
wire cdxi2707m = reg_0_3&cdxi1751m;
wire cdxi2708m = reg_0_3&cdxi1752m;
wire cdxi2709m = reg_0_3&cdxi1753m;
wire cdxi2710m = reg_0_6&cdxi1646m;
wire cdxi2711m = reg_0_5&cdxi1680m;
wire cdxi2712m = reg_0_5&cdxi1681m;
wire cdxi2713m = reg_0_4&cdxi1576m;
wire cdxi2714m = reg_0_4&cdxi1577m;
wire cdxi2715m = reg_0_4&cdxi1578m;
wire cdxi2716m = reg_0_3&cdxi1754m;
wire cdxi2717m = reg_0_3&cdxi1755m;
wire cdxi2718m = reg_0_3&cdxi1756m;
wire cdxi2719m = reg_0_3&cdxi1757m;
wire cdxi2720m = reg_0_7&cdxi1703m;
wire cdxi2721m = reg_0_6&cdxi1635m;
wire cdxi2722m = reg_0_5&cdxi1669m;
wire cdxi2723m = reg_0_4&cdxi1565m;
wire cdxi2724m = reg_0_3&cdxi1743m;
wire cdxi2725m = (cdxi2695m ^ cdxi2696m ^ cdxi2697m ^ cdxi2698m ^ cdxi2699m ^ cdxi2700m ^ cdxi2701m ^ cdxi2702m ^ cdxi2703m ^ cdxi2704m ^ cdxi2705m ^ cdxi2706m ^ cdxi2707m ^ cdxi2708m ^ cdxi2709m ^ cdxi2710m ^ cdxi2711m ^ cdxi2712m ^ cdxi2713m ^ cdxi2714m ^ cdxi2715m ^ cdxi2716m ^ cdxi2717m ^ cdxi2718m ^ cdxi2719m ^ cdxi2720m ^ cdxi2721m ^ cdxi2722m ^ cdxi2723m ^ cdxi2724m ^ cdxi2694m);
wire cdxi2726m = reg_0_0&cdxi2725m;
wire cdxi2727m = cdxi185m&cdxi2491m;
wire cdxi2728m = reg_0_1&cdxi2524m;
wire cdxi2729m = cdxi185m&cdxi2559m;
wire cdxi2730m = reg_0_1&cdxi2592m;
wire cdxi2731m = cdxi361m&cdxi1548m ^ r116m;
wire cdxi2732m = cdxi1374m&cdxi271m;
wire cdxi2733m = cdxi1013m&cdxi230m;
wire cdxi2734m = cdxi361m&cdxi658m;
wire cdxi2735m = cdxi361m&cdxi659m;
wire cdxi2736m = cdxi361m&cdxi660m;
wire cdxi2737m = cdxi1548m&r13m;
wire cdxi2738m = cdxi601m&cdxi737m;
wire cdxi2739m = cdxi1160m&r16m;
wire cdxi2740m = cdxi1374m&r17m;
wire cdxi2741m = cdxi384m&cdxi623m;
wire cdxi2742m = cdxi1410m&r20m;
wire cdxi2743m = cdxi1013m&r21m;
wire cdxi2744m = cdxi361m&cdxi661m;
wire cdxi2745m = cdxi361m&cdxi662m;
wire cdxi2746m = cdxi361m&cdxi663m;
wire cdxi2747m = cdxi657m&r44m;
wire cdxi2748m = cdxi485m&r45m;
wire cdxi2749m = cdxi638m&r46m;
wire cdxi2750m = cdxi425m&r50m;
wire cdxi2751m = cdxi601m&r51m;
wire cdxi2752m = cdxi582m&r52m;
wire cdxi2753m = cdxi563m&r56m;
wire cdxi2754m = cdxi384m&r57m;
wire cdxi2755m = cdxi524m&r58m;
wire cdxi2756m = cdxi361m&r62m;
wire cdxi2757m = cdxi207m&r86m;
wire cdxi2758m = cdxi218m&r87m;
wire cdxi2759m = cdxi240m&r88m;
wire cdxi2760m = cdxi184m&r92m;
wire cdxi2761m = cdxi219m&r96m;
wire cdxi2762m = (cdxi2731m ^ cdxi2732m ^ cdxi2733m ^ cdxi2734m ^ cdxi2735m ^ cdxi2736m ^ cdxi2737m ^ cdxi2738m ^ cdxi2739m ^ cdxi2740m ^ cdxi2741m ^ cdxi2742m ^ cdxi2743m ^ cdxi2744m ^ cdxi2745m ^ cdxi2746m ^ cdxi2747m ^ cdxi2748m ^ cdxi2749m ^ cdxi2750m ^ cdxi2751m ^ cdxi2752m ^ cdxi2753m ^ cdxi2754m ^ cdxi2755m ^ cdxi2756m ^ cdxi2757m ^ cdxi2758m ^ cdxi2759m ^ cdxi2760m ^ cdxi2761m);
wire cdxi2763m = cdxi185m&cdxi2762m;
wire cdxi2764m = (reg_0_124);
wire cdxi2765m = reg_0_3&reg_0_5&reg_0_6&cdxi276m;
wire cdxi2766m = reg_0_2&cdxi1566m;
wire cdxi2767m = reg_0_2&cdxi1567m;
wire cdxi2768m = reg_0_2&cdxi1568m;
wire cdxi2769m = reg_0_2&cdxi1569m;
wire cdxi2770m = reg_0_5&cdxi1466m;
wire cdxi2771m = reg_0_3&reg_0_6&cdxi746m;
wire cdxi2772m = reg_0_3&reg_0_5&reg_0_7&cdxi224m;
wire cdxi2773m = reg_0_3&reg_0_5&reg_0_6&cdxi275m;
wire cdxi2774m = reg_0_2&cdxi1570m;
wire cdxi2775m = reg_0_2&cdxi1571m;
wire cdxi2776m = reg_0_2&cdxi1572m;
wire cdxi2777m = reg_0_2&cdxi1573m;
wire cdxi2778m = reg_0_2&cdxi1574m;
wire cdxi2779m = reg_0_2&cdxi1575m;
wire cdxi2780m = reg_0_6&cdxi1438m;
wire cdxi2781m = reg_0_5&cdxi1472m;
wire cdxi2782m = reg_0_5&cdxi1473m;
wire cdxi2783m = reg_0_3&reg_0_7&cdxi724m;
wire cdxi2784m = reg_0_3&reg_0_6&cdxi742m;
wire cdxi2785m = reg_0_3&reg_0_5&cdxi1069m;
wire cdxi2786m = reg_0_2&cdxi1576m;
wire cdxi2787m = reg_0_2&cdxi1577m;
wire cdxi2788m = reg_0_2&cdxi1578m;
wire cdxi2789m = reg_0_2&cdxi1579m;
wire cdxi2790m = reg_0_7&cdxi1392m;
wire cdxi2791m = reg_0_6&cdxi1427m;
wire cdxi2792m = reg_0_5&cdxi1461m;
wire cdxi2793m = reg_0_3&cdxi2221m;
wire cdxi2794m = reg_0_2&cdxi1565m;
wire cdxi2795m = (cdxi2765m ^ cdxi2766m ^ cdxi2767m ^ cdxi2768m ^ cdxi2769m ^ cdxi2770m ^ cdxi2771m ^ cdxi2772m ^ cdxi2773m ^ cdxi2774m ^ cdxi2775m ^ cdxi2776m ^ cdxi2777m ^ cdxi2778m ^ cdxi2779m ^ cdxi2780m ^ cdxi2781m ^ cdxi2782m ^ cdxi2783m ^ cdxi2784m ^ cdxi2785m ^ cdxi2786m ^ cdxi2787m ^ cdxi2788m ^ cdxi2789m ^ cdxi2790m ^ cdxi2791m ^ cdxi2792m ^ cdxi2793m ^ cdxi2794m ^ cdxi2764m);
wire cdxi2796m = reg_0_1&cdxi2795m;
wire cdxi2797m = cdxi185m&cdxi2692m;
wire cdxi2798m = reg_0_1&cdxi2725m;
wire cdxi2799m = cdxi825m&cdxi1268m ^ r121m;
wire cdxi2800m = cdxi361m&cdxi1268m;
wire cdxi2801m = cdxi362m&cdxi1268m;
wire cdxi2802m = cdxi363m&cdxi1268m;
wire cdxi2803m = cdxi825m&cdxi657m;
wire cdxi2804m = cdxi825m&cdxi562m;
wire cdxi2805m = cdxi825m&cdxi466m;
wire cdxi2806m = cdxi362m&cdxi657m;
wire cdxi2807m = cdxi361m&cdxi1269m;
wire cdxi2808m = cdxi1835m&cdxi271m;
wire cdxi2809m = cdxi363m&cdxi1653m;
wire cdxi2810m = cdxi825m&cdxi758m;
wire cdxi2811m = cdxi825m&cdxi759m;
wire cdxi2812m = cdxi825m&cdxi760m;
wire cdxi2813m = cdxi405m&cdxi1056m;
wire cdxi2814m = cdxi977m&cdxi430m;
wire cdxi2815m = cdxi361m&cdxi1273m;
wire cdxi2816m = cdxi361m&cdxi1274m;
wire cdxi2817m = cdxi361m&cdxi1275m;
wire cdxi2818m = cdxi406m&cdxi1449m;
wire cdxi2819m = cdxi901m&cdxi567m;
wire cdxi2820m = cdxi2325m&r16m;
wire cdxi2821m = cdxi1835m&r17m;
wire cdxi2822m = cdxi363m&cdxi1657m;
wire cdxi2823m = cdxi363m&cdxi1658m;
wire cdxi2824m = cdxi363m&cdxi1659m;
wire cdxi2825m = cdxi825m&cdxi761m;
wire cdxi2826m = cdxi825m&cdxi762m;
wire cdxi2827m = cdxi825m&cdxi763m;
wire cdxi2828m = cdxi466m&cdxi951m;
wire cdxi2829m = cdxi1196m&r29m;
wire cdxi2830m = cdxi405m&cdxi1062m;
wire cdxi2831m = cdxi405m&cdxi1063m;
wire cdxi2832m = cdxi1050m&r33m;
wire cdxi2833m = cdxi504m&cdxi1207m;
wire cdxi2834m = cdxi977m&r36m;
wire cdxi2835m = cdxi938m&r38m;
wire cdxi2836m = cdxi900m&r39m;
wire cdxi2837m = cdxi822m&r42m;
wire cdxi2838m = cdxi1051m&r43m;
wire cdxi2839m = cdxi1124m&r45m;
wire cdxi2840m = cdxi978m&r46m;
wire cdxi2841m = cdxi939m&r48m;
wire cdxi2842m = cdxi901m&r49m;
wire cdxi2843m = cdxi823m&r52m;
wire cdxi2844m = cdxi940m&r54m;
wire cdxi2845m = cdxi902m&r55m;
wire cdxi2846m = cdxi824m&r58m;
wire cdxi2847m = cdxi825m&r61m;
wire cdxi2848m = cdxi657m&r63m;
wire cdxi2849m = cdxi562m&r65m;
wire cdxi2850m = cdxi466m&r66m;
wire cdxi2851m = cdxi425m&r68m;
wire cdxi2852m = cdxi601m&r69m;
wire cdxi2853m = cdxi405m&r72m;
wire cdxi2854m = cdxi563m&r74m;
wire cdxi2855m = cdxi384m&r75m;
wire cdxi2856m = cdxi504m&r78m;
wire cdxi2857m = cdxi361m&r81m;
wire cdxi2858m = cdxi426m&r84m;
wire cdxi2859m = cdxi385m&r85m;
wire cdxi2860m = cdxi406m&r88m;
wire cdxi2861m = cdxi362m&r91m;
wire cdxi2862m = cdxi363m&r95m;
wire cdxi2863m = cdxi207m&r99m;
wire cdxi2864m = cdxi218m&r100m;
wire cdxi2865m = cdxi196m&r103m;
wire cdxi2866m = cdxi184m&r106m;
wire cdxi2867m = cdxi219m&r110m;
wire cdxi2868m = cdxi185m&r115m;
wire cdxi2869m = (cdxi2799m ^ cdxi2807m ^ cdxi2808m ^ cdxi2809m ^ cdxi2810m ^ cdxi2811m ^ cdxi2812m ^ cdxi2813m ^ cdxi2814m ^ cdxi2815m ^ cdxi2816m ^ cdxi2817m ^ cdxi2818m ^ cdxi2819m ^ cdxi2820m ^ cdxi2821m ^ cdxi2822m ^ cdxi2823m ^ cdxi2824m ^ cdxi2825m ^ cdxi2826m ^ cdxi2827m ^ cdxi2828m ^ cdxi2829m ^ cdxi2830m ^ cdxi2831m ^ cdxi2832m ^ cdxi2833m ^ cdxi2834m ^ cdxi2835m ^ cdxi2836m ^ cdxi2837m ^ cdxi2838m ^ cdxi2839m ^ cdxi2840m ^ cdxi2841m ^ cdxi2842m ^ cdxi2843m ^ cdxi2844m ^ cdxi2845m ^ cdxi2846m ^ cdxi2847m ^ cdxi2848m ^ cdxi2849m ^ cdxi2850m ^ cdxi2851m ^ cdxi2852m ^ cdxi2853m ^ cdxi2854m ^ cdxi2855m ^ cdxi2856m ^ cdxi2857m ^ cdxi2858m ^ cdxi2859m ^ cdxi2860m ^ cdxi2861m ^ cdxi2862m ^ cdxi2863m ^ cdxi2864m ^ cdxi2865m ^ cdxi2866m ^ cdxi2867m ^ cdxi2868m);
wire cdxi2870m = a0&cdxi2869m;
wire cdxi2871m = (reg_0_108);
wire cdxi2872m = (reg_0_111);
wire cdxi2873m = (reg_0_118);
wire cdxi2874m = (reg_0_129);
wire cdxi2875m = reg_0_2&reg_0_3&cdxi1286m;
wire cdxi2876m = reg_0_1&cdxi2562m;
wire cdxi2877m = reg_0_1&cdxi2563m;
wire cdxi2878m = reg_0_1&cdxi2564m;
wire cdxi2879m = reg_0_1&cdxi2565m;
wire cdxi2880m = reg_0_1&cdxi2566m;
wire cdxi2881m = reg_0_3&cdxi2158m;
wire cdxi2882m = reg_0_2&reg_0_4&cdxi1219m;
wire cdxi2883m = reg_0_2&reg_0_3&cdxi1290m;
wire cdxi2884m = reg_0_2&reg_0_3&cdxi1291m;
wire cdxi2885m = reg_0_2&reg_0_3&cdxi1292m;
wire cdxi2886m = reg_0_1&cdxi2567m;
wire cdxi2887m = reg_0_1&cdxi2568m;
wire cdxi2888m = reg_0_1&cdxi2569m;
wire cdxi2889m = reg_0_1&cdxi2570m;
wire cdxi2890m = reg_0_1&cdxi2571m;
wire cdxi2891m = reg_0_1&cdxi2572m;
wire cdxi2892m = reg_0_1&cdxi2573m;
wire cdxi2893m = reg_0_1&cdxi2574m;
wire cdxi2894m = reg_0_1&cdxi2575m;
wire cdxi2895m = reg_0_1&cdxi2576m;
wire cdxi2896m = reg_0_4&reg_0_6&cdxi970m;
wire cdxi2897m = reg_0_3&cdxi2168m;
wire cdxi2898m = reg_0_3&cdxi2169m;
wire cdxi2899m = reg_0_3&cdxi2170m;
wire cdxi2900m = reg_0_2&reg_0_6&cdxi1153m;
wire cdxi2901m = reg_0_2&reg_0_4&cdxi1225m;
wire cdxi2902m = reg_0_2&reg_0_4&cdxi1226m;
wire cdxi2903m = reg_0_2&reg_0_3&cdxi1296m;
wire cdxi2904m = reg_0_2&reg_0_3&cdxi1297m;
wire cdxi2905m = reg_0_2&reg_0_3&cdxi1298m;
wire cdxi2906m = reg_0_1&cdxi2577m;
wire cdxi2907m = reg_0_1&cdxi2578m;
wire cdxi2908m = reg_0_1&cdxi2579m;
wire cdxi2909m = reg_0_1&cdxi2580m;
wire cdxi2910m = reg_0_1&cdxi2581m;
wire cdxi2911m = reg_0_1&cdxi2582m;
wire cdxi2912m = reg_0_1&cdxi2583m;
wire cdxi2913m = reg_0_1&cdxi2584m;
wire cdxi2914m = reg_0_1&cdxi2585m;
wire cdxi2915m = reg_0_1&cdxi2586m;
wire cdxi2916m = reg_0_6&reg_0_7&cdxi843m;
wire cdxi2917m = reg_0_4&reg_0_7&cdxi920m;
wire cdxi2918m = reg_0_4&reg_0_6&cdxi959m;
wire cdxi2919m = reg_0_3&cdxi2178m;
wire cdxi2920m = reg_0_3&cdxi2179m;
wire cdxi2921m = reg_0_3&cdxi2180m;
wire cdxi2922m = reg_0_2&reg_0_7&cdxi1105m;
wire cdxi2923m = reg_0_2&reg_0_6&cdxi1142m;
wire cdxi2924m = reg_0_2&reg_0_4&cdxi1214m;
wire cdxi2925m = reg_0_2&reg_0_3&cdxi1285m;
wire cdxi2926m = reg_0_1&cdxi2587m;
wire cdxi2927m = reg_0_1&cdxi2588m;
wire cdxi2928m = reg_0_1&cdxi2589m;
wire cdxi2929m = reg_0_1&cdxi2590m;
wire cdxi2930m = reg_0_1&cdxi2591m;
wire cdxi2931m = reg_0_7&cdxi1870m;
wire cdxi2932m = reg_0_6&cdxi2871m;
wire cdxi2933m = reg_0_4&cdxi2872m;
wire cdxi2934m = reg_0_3&cdxi2152m;
wire cdxi2935m = reg_0_2&cdxi2873m;
wire cdxi2936m = reg_0_1&cdxi2561m;
wire cdxi2937m = (cdxi2875m ^ cdxi2876m ^ cdxi2877m ^ cdxi2878m ^ cdxi2879m ^ cdxi2880m ^ cdxi2881m ^ cdxi2882m ^ cdxi2883m ^ cdxi2884m ^ cdxi2885m ^ cdxi2886m ^ cdxi2887m ^ cdxi2888m ^ cdxi2889m ^ cdxi2890m ^ cdxi2891m ^ cdxi2892m ^ cdxi2893m ^ cdxi2894m ^ cdxi2895m ^ cdxi2896m ^ cdxi2897m ^ cdxi2898m ^ cdxi2899m ^ cdxi2900m ^ cdxi2901m ^ cdxi2902m ^ cdxi2903m ^ cdxi2904m ^ cdxi2905m ^ cdxi2906m ^ cdxi2907m ^ cdxi2908m ^ cdxi2909m ^ cdxi2910m ^ cdxi2911m ^ cdxi2912m ^ cdxi2913m ^ cdxi2914m ^ cdxi2915m ^ cdxi2916m ^ cdxi2917m ^ cdxi2918m ^ cdxi2919m ^ cdxi2920m ^ cdxi2921m ^ cdxi2922m ^ cdxi2923m ^ cdxi2924m ^ cdxi2925m ^ cdxi2926m ^ cdxi2927m ^ cdxi2928m ^ cdxi2929m ^ cdxi2930m ^ cdxi2931m ^ cdxi2932m ^ cdxi2933m ^ cdxi2934m ^ cdxi2935m ^ cdxi2936m ^ cdxi2874m);
wire cdxi2938m = reg_0_0&cdxi2937m;
wire cdxi2939m = cdxi825m&cdxi1548m ^ r122m;
wire cdxi2940m = cdxi361m&cdxi1548m;
wire cdxi2941m = cdxi362m&cdxi1548m;
wire cdxi2942m = cdxi363m&cdxi1548m;
wire cdxi2943m = cdxi825m&cdxi485m;
wire cdxi2944m = cdxi825m&cdxi638m;
wire cdxi2945m = cdxi1904m&cdxi208m;
wire cdxi2946m = cdxi1905m&cdxi271m;
wire cdxi2947m = cdxi363m&cdxi1549m;
wire cdxi2948m = cdxi825m&cdxi658m;
wire cdxi2949m = cdxi825m&cdxi659m;
wire cdxi2950m = cdxi825m&cdxi660m;
wire cdxi2951m = cdxi582m&cdxi1056m;
wire cdxi2952m = cdxi1013m&cdxi430m;
wire cdxi2953m = cdxi900m&cdxi489m;
wire cdxi2954m = cdxi1974m&r11m;
wire cdxi2955m = cdxi1904m&r12m;
wire cdxi2956m = cdxi446m&cdxi1449m;
wire cdxi2957m = cdxi2806m&r15m;
wire cdxi2958m = cdxi1975m&r16m;
wire cdxi2959m = cdxi1905m&r17m;
wire cdxi2960m = cdxi902m&cdxi623m;
wire cdxi2961m = cdxi363m&cdxi1554m;
wire cdxi2962m = cdxi363m&cdxi1555m;
wire cdxi2963m = cdxi825m&cdxi661m;
wire cdxi2964m = cdxi825m&cdxi662m;
wire cdxi2965m = cdxi825m&cdxi663m;
wire cdxi2966m = cdxi638m&cdxi951m;
wire cdxi2967m = cdxi1196m&r30m;
wire cdxi2968m = cdxi1160m&r31m;
wire cdxi2969m = cdxi582m&cdxi1063m;
wire cdxi2970m = cdxi1050m&r34m;
wire cdxi2971m = cdxi1410m&r35m;
wire cdxi2972m = cdxi1013m&r36m;
wire cdxi2973m = cdxi938m&r40m;
wire cdxi2974m = cdxi900m&r41m;
wire cdxi2975m = cdxi861m&r42m;
wire cdxi2976m = cdxi1051m&r44m;
wire cdxi2977m = cdxi1161m&r45m;
wire cdxi2978m = cdxi1014m&r46m;
wire cdxi2979m = cdxi939m&r50m;
wire cdxi2980m = cdxi901m&r51m;
wire cdxi2981m = cdxi862m&r52m;
wire cdxi2982m = cdxi940m&r56m;
wire cdxi2983m = cdxi902m&r57m;
wire cdxi2984m = cdxi863m&r58m;
wire cdxi2985m = cdxi825m&r62m;
wire cdxi2986m = cdxi657m&r64m;
wire cdxi2987m = cdxi485m&r65m;
wire cdxi2988m = cdxi638m&r66m;
wire cdxi2989m = cdxi425m&r70m;
wire cdxi2990m = cdxi601m&r71m;
wire cdxi2991m = cdxi582m&r72m;
wire cdxi2992m = cdxi563m&r76m;
wire cdxi2993m = cdxi384m&r77m;
wire cdxi2994m = cdxi524m&r78m;
wire cdxi2995m = cdxi361m&r82m;
wire cdxi2996m = cdxi426m&r86m;
wire cdxi2997m = cdxi385m&r87m;
wire cdxi2998m = cdxi446m&r88m;
wire cdxi2999m = cdxi362m&r92m;
wire cdxi3000m = cdxi363m&r96m;
wire cdxi3001m = cdxi207m&r101m;
wire cdxi3002m = cdxi218m&r102m;
wire cdxi3003m = cdxi240m&r103m;
wire cdxi3004m = cdxi184m&r107m;
wire cdxi3005m = cdxi219m&r111m;
wire cdxi3006m = cdxi185m&r116m;
wire cdxi3007m = (cdxi2939m ^ cdxi2945m ^ cdxi2946m ^ cdxi2947m ^ cdxi2948m ^ cdxi2949m ^ cdxi2950m ^ cdxi2951m ^ cdxi2952m ^ cdxi2953m ^ cdxi2954m ^ cdxi2955m ^ cdxi2956m ^ cdxi2957m ^ cdxi2958m ^ cdxi2959m ^ cdxi2960m ^ cdxi2961m ^ cdxi2962m ^ cdxi2963m ^ cdxi2964m ^ cdxi2965m ^ cdxi2966m ^ cdxi2967m ^ cdxi2968m ^ cdxi2969m ^ cdxi2970m ^ cdxi2971m ^ cdxi2972m ^ cdxi2973m ^ cdxi2974m ^ cdxi2975m ^ cdxi2976m ^ cdxi2977m ^ cdxi2978m ^ cdxi2979m ^ cdxi2980m ^ cdxi2981m ^ cdxi2982m ^ cdxi2983m ^ cdxi2984m ^ cdxi2985m ^ cdxi2986m ^ cdxi2987m ^ cdxi2988m ^ cdxi2989m ^ cdxi2990m ^ cdxi2991m ^ cdxi2992m ^ cdxi2993m ^ cdxi2994m ^ cdxi2995m ^ cdxi2996m ^ cdxi2997m ^ cdxi2998m ^ cdxi2999m ^ cdxi3000m ^ cdxi3001m ^ cdxi3002m ^ cdxi3003m ^ cdxi3004m ^ cdxi3005m ^ cdxi3006m);
wire cdxi3008m = a0&cdxi3007m;
wire cdxi3009m = (reg_0_119);
wire cdxi3010m = (reg_0_130);
wire cdxi3011m = reg_0_2&reg_0_3&reg_0_5&reg_0_6&cdxi213m;
wire cdxi3012m = reg_0_1&cdxi2765m;
wire cdxi3013m = reg_0_1&cdxi2766m;
wire cdxi3014m = reg_0_1&cdxi2767m;
wire cdxi3015m = reg_0_1&cdxi2768m;
wire cdxi3016m = reg_0_1&cdxi2769m;
wire cdxi3017m = reg_0_3&cdxi2228m;
wire cdxi3018m = reg_0_2&reg_0_5&cdxi1219m;
wire cdxi3019m = reg_0_2&reg_0_3&reg_0_6&cdxi498m;
wire cdxi3020m = reg_0_2&reg_0_3&reg_0_5&reg_0_7&cdxi394m;
wire cdxi3021m = reg_0_2&reg_0_3&reg_0_5&reg_0_6&cdxi212m;
wire cdxi3022m = reg_0_1&cdxi2770m;
wire cdxi3023m = reg_0_1&cdxi2771m;
wire cdxi3024m = reg_0_1&cdxi2772m;
wire cdxi3025m = reg_0_1&cdxi2773m;
wire cdxi3026m = reg_0_1&cdxi2774m;
wire cdxi3027m = reg_0_1&cdxi2775m;
wire cdxi3028m = reg_0_1&cdxi2776m;
wire cdxi3029m = reg_0_1&cdxi2777m;
wire cdxi3030m = reg_0_1&cdxi2778m;
wire cdxi3031m = reg_0_1&cdxi2779m;
wire cdxi3032m = reg_0_5&reg_0_6&cdxi970m;
wire cdxi3033m = reg_0_3&cdxi2238m;
wire cdxi3034m = reg_0_3&cdxi2239m;
wire cdxi3035m = reg_0_3&cdxi2240m;
wire cdxi3036m = reg_0_2&reg_0_6&cdxi1189m;
wire cdxi3037m = reg_0_2&reg_0_5&cdxi1225m;
wire cdxi3038m = reg_0_2&reg_0_5&cdxi1226m;
wire cdxi3039m = reg_0_2&reg_0_3&reg_0_7&cdxi1031m;
wire cdxi3040m = reg_0_2&reg_0_3&reg_0_6&cdxi494m;
wire cdxi3041m = reg_0_2&reg_0_3&reg_0_5&cdxi1068m;
wire cdxi3042m = reg_0_1&cdxi2780m;
wire cdxi3043m = reg_0_1&cdxi2781m;
wire cdxi3044m = reg_0_1&cdxi2782m;
wire cdxi3045m = reg_0_1&cdxi2783m;
wire cdxi3046m = reg_0_1&cdxi2784m;
wire cdxi3047m = reg_0_1&cdxi2785m;
wire cdxi3048m = reg_0_1&cdxi2786m;
wire cdxi3049m = reg_0_1&cdxi2787m;
wire cdxi3050m = reg_0_1&cdxi2788m;
wire cdxi3051m = reg_0_1&cdxi2789m;
wire cdxi3052m = reg_0_6&cdxi2037m;
wire cdxi3053m = reg_0_5&reg_0_7&cdxi920m;
wire cdxi3054m = reg_0_5&reg_0_6&cdxi959m;
wire cdxi3055m = reg_0_3&cdxi2248m;
wire cdxi3056m = reg_0_3&cdxi2249m;
wire cdxi3057m = reg_0_3&cdxi2250m;
wire cdxi3058m = reg_0_2&reg_0_7&cdxi1939m;
wire cdxi3059m = reg_0_2&reg_0_6&cdxi1178m;
wire cdxi3060m = reg_0_2&reg_0_5&cdxi1214m;
wire cdxi3061m = reg_0_2&reg_0_3&cdxi2220m;
wire cdxi3062m = reg_0_1&cdxi2790m;
wire cdxi3063m = reg_0_1&cdxi2791m;
wire cdxi3064m = reg_0_1&cdxi2792m;
wire cdxi3065m = reg_0_1&cdxi2793m;
wire cdxi3066m = reg_0_1&cdxi2794m;
wire cdxi3067m = reg_0_7&cdxi1940m;
wire cdxi3068m = reg_0_6&cdxi2011m;
wire cdxi3069m = reg_0_5&cdxi2872m;
wire cdxi3070m = reg_0_3&cdxi2222m;
wire cdxi3071m = reg_0_2&cdxi3009m;
wire cdxi3072m = reg_0_1&cdxi2764m;
wire cdxi3073m = (cdxi3011m ^ cdxi3012m ^ cdxi3013m ^ cdxi3014m ^ cdxi3015m ^ cdxi3016m ^ cdxi3017m ^ cdxi3018m ^ cdxi3019m ^ cdxi3020m ^ cdxi3021m ^ cdxi3022m ^ cdxi3023m ^ cdxi3024m ^ cdxi3025m ^ cdxi3026m ^ cdxi3027m ^ cdxi3028m ^ cdxi3029m ^ cdxi3030m ^ cdxi3031m ^ cdxi3032m ^ cdxi3033m ^ cdxi3034m ^ cdxi3035m ^ cdxi3036m ^ cdxi3037m ^ cdxi3038m ^ cdxi3039m ^ cdxi3040m ^ cdxi3041m ^ cdxi3042m ^ cdxi3043m ^ cdxi3044m ^ cdxi3045m ^ cdxi3046m ^ cdxi3047m ^ cdxi3048m ^ cdxi3049m ^ cdxi3050m ^ cdxi3051m ^ cdxi3052m ^ cdxi3053m ^ cdxi3054m ^ cdxi3055m ^ cdxi3056m ^ cdxi3057m ^ cdxi3058m ^ cdxi3059m ^ cdxi3060m ^ cdxi3061m ^ cdxi3062m ^ cdxi3063m ^ cdxi3064m ^ cdxi3065m ^ cdxi3066m ^ cdxi3067m ^ cdxi3068m ^ cdxi3069m ^ cdxi3070m ^ cdxi3071m ^ cdxi3072m ^ cdxi3010m);
wire cdxi3074m = reg_0_0&cdxi3073m;
wire cdxi3075m = cdxi1763m&cdxi657m ^ r123m;
wire cdxi3076m = cdxi1304m&cdxi657m;
wire cdxi3077m = cdxi406m&cdxi1548m;
wire cdxi3078m = cdxi363m&cdxi1232m;
wire cdxi3079m = cdxi363m&cdxi1479m;
wire cdxi3080m = cdxi2045m&cdxi208m;
wire cdxi3081m = cdxi2046m&cdxi271m;
wire cdxi3082m = cdxi363m&cdxi1727m;
wire cdxi3083m = cdxi363m&cdxi1728m;
wire cdxi3084m = cdxi363m&cdxi1729m;
wire cdxi3085m = cdxi363m&cdxi1730m;
wire cdxi3086m = cdxi445m&cdxi1056m;
wire cdxi3087m = cdxi524m&cdxi1273m;
wire cdxi3088m = cdxi977m&cdxi489m;
wire cdxi3089m = cdxi219m&cdxi2400m;
wire cdxi3090m = cdxi2045m&r12m;
wire cdxi3091m = cdxi1014m&cdxi567m;
wire cdxi3092m = cdxi2115m&r15m;
wire cdxi3093m = cdxi2324m&r16m;
wire cdxi3094m = cdxi2046m&r17m;
wire cdxi3095m = cdxi363m&cdxi1731m;
wire cdxi3096m = cdxi363m&cdxi1732m;
wire cdxi3097m = cdxi363m&cdxi1733m;
wire cdxi3098m = cdxi363m&cdxi1734m;
wire cdxi3099m = cdxi363m&cdxi1735m;
wire cdxi3100m = cdxi363m&cdxi1736m;
wire cdxi3101m = cdxi1548m&r29m;
wire cdxi3102m = cdxi1268m&r30m;
wire cdxi3103m = cdxi445m&cdxi1062m;
wire cdxi3104m = cdxi445m&cdxi1063m;
wire cdxi3105m = cdxi1050m&r37m;
wire cdxi3106m = cdxi1410m&r38m;
wire cdxi3107m = cdxi1013m&r39m;
wire cdxi3108m = cdxi1339m&r40m;
wire cdxi3109m = cdxi977m&r41m;
wire cdxi3110m = cdxi1304m&r42m;
wire cdxi3111m = cdxi1051m&r47m;
wire cdxi3112m = cdxi1161m&r48m;
wire cdxi3113m = cdxi1014m&r49m;
wire cdxi3114m = cdxi1124m&r50m;
wire cdxi3115m = cdxi978m&r51m;
wire cdxi3116m = cdxi1233m&r52m;
wire cdxi3117m = cdxi940m&r59m;
wire cdxi3118m = cdxi902m&r60m;
wire cdxi3119m = cdxi863m&r61m;
wire cdxi3120m = cdxi824m&r62m;
wire cdxi3121m = cdxi657m&r67m;
wire cdxi3122m = cdxi485m&r68m;
wire cdxi3123m = cdxi638m&r69m;
wire cdxi3124m = cdxi562m&r70m;
wire cdxi3125m = cdxi466m&r71m;
wire cdxi3126m = cdxi445m&r72m;
wire cdxi3127m = cdxi563m&r79m;
wire cdxi3128m = cdxi384m&r80m;
wire cdxi3129m = cdxi524m&r81m;
wire cdxi3130m = cdxi504m&r82m;
wire cdxi3131m = cdxi426m&r89m;
wire cdxi3132m = cdxi385m&r90m;
wire cdxi3133m = cdxi446m&r91m;
wire cdxi3134m = cdxi406m&r92m;
wire cdxi3135m = cdxi363m&r97m;
wire cdxi3136m = cdxi207m&r104m;
wire cdxi3137m = cdxi218m&r105m;
wire cdxi3138m = cdxi240m&r106m;
wire cdxi3139m = cdxi196m&r107m;
wire cdxi3140m = cdxi219m&r112m;
wire cdxi3141m = cdxi185m&r117m;
wire cdxi3142m = (cdxi3075m ^ cdxi3080m ^ cdxi3081m ^ cdxi3082m ^ cdxi3083m ^ cdxi3084m ^ cdxi3085m ^ cdxi3086m ^ cdxi3087m ^ cdxi3088m ^ cdxi3089m ^ cdxi3090m ^ cdxi3091m ^ cdxi3092m ^ cdxi3093m ^ cdxi3094m ^ cdxi3095m ^ cdxi3096m ^ cdxi3097m ^ cdxi3098m ^ cdxi3099m ^ cdxi3100m ^ cdxi3101m ^ cdxi3102m ^ cdxi3103m ^ cdxi3104m ^ cdxi3105m ^ cdxi3106m ^ cdxi3107m ^ cdxi3108m ^ cdxi3109m ^ cdxi3110m ^ cdxi3111m ^ cdxi3112m ^ cdxi3113m ^ cdxi3114m ^ cdxi3115m ^ cdxi3116m ^ cdxi3117m ^ cdxi3118m ^ cdxi3119m ^ cdxi3120m ^ cdxi3121m ^ cdxi3122m ^ cdxi3123m ^ cdxi3124m ^ cdxi3125m ^ cdxi3126m ^ cdxi3127m ^ cdxi3128m ^ cdxi3129m ^ cdxi3130m ^ cdxi3131m ^ cdxi3132m ^ cdxi3133m ^ cdxi3134m ^ cdxi3135m ^ cdxi3136m ^ cdxi3137m ^ cdxi3138m ^ cdxi3139m ^ cdxi3140m ^ cdxi3141m);
wire cdxi3143m = a0&cdxi3142m;
wire cdxi3144m = (reg_0_113);
wire cdxi3145m = (reg_0_131);
wire cdxi3146m = reg_0_2&cdxi2426m;
wire cdxi3147m = reg_0_1&cdxi2628m;
wire cdxi3148m = reg_0_1&cdxi2629m;
wire cdxi3149m = reg_0_1&cdxi2630m;
wire cdxi3150m = reg_0_1&cdxi2631m;
wire cdxi3151m = reg_0_1&cdxi2632m;
wire cdxi3152m = reg_0_4&cdxi2228m;
wire cdxi3153m = reg_0_2&cdxi2431m;
wire cdxi3154m = reg_0_2&cdxi2432m;
wire cdxi3155m = reg_0_2&cdxi2433m;
wire cdxi3156m = reg_0_2&cdxi2434m;
wire cdxi3157m = reg_0_1&cdxi2633m;
wire cdxi3158m = reg_0_1&cdxi2634m;
wire cdxi3159m = reg_0_1&cdxi2635m;
wire cdxi3160m = reg_0_1&cdxi2636m;
wire cdxi3161m = reg_0_1&cdxi2637m;
wire cdxi3162m = reg_0_1&cdxi2638m;
wire cdxi3163m = reg_0_1&cdxi2639m;
wire cdxi3164m = reg_0_1&cdxi2640m;
wire cdxi3165m = reg_0_1&cdxi2641m;
wire cdxi3166m = reg_0_1&cdxi2642m;
wire cdxi3167m = reg_0_5&cdxi2168m;
wire cdxi3168m = reg_0_4&cdxi2238m;
wire cdxi3169m = reg_0_4&cdxi2239m;
wire cdxi3170m = reg_0_4&cdxi2240m;
wire cdxi3171m = reg_0_2&cdxi2441m;
wire cdxi3172m = reg_0_2&cdxi2442m;
wire cdxi3173m = reg_0_2&cdxi2443m;
wire cdxi3174m = reg_0_2&cdxi2444m;
wire cdxi3175m = reg_0_2&cdxi2445m;
wire cdxi3176m = reg_0_2&cdxi2446m;
wire cdxi3177m = reg_0_1&cdxi2643m;
wire cdxi3178m = reg_0_1&cdxi2644m;
wire cdxi3179m = reg_0_1&cdxi2645m;
wire cdxi3180m = reg_0_1&cdxi2646m;
wire cdxi3181m = reg_0_1&cdxi2647m;
wire cdxi3182m = reg_0_1&cdxi2648m;
wire cdxi3183m = reg_0_1&cdxi2649m;
wire cdxi3184m = reg_0_1&cdxi2650m;
wire cdxi3185m = reg_0_1&cdxi2651m;
wire cdxi3186m = reg_0_1&cdxi2652m;
wire cdxi3187m = reg_0_6&reg_0_7&cdxi1798m;
wire cdxi3188m = reg_0_5&cdxi2178m;
wire cdxi3189m = reg_0_5&cdxi2179m;
wire cdxi3190m = reg_0_4&cdxi2248m;
wire cdxi3191m = reg_0_4&cdxi2249m;
wire cdxi3192m = reg_0_4&cdxi2250m;
wire cdxi3193m = reg_0_2&cdxi2451m;
wire cdxi3194m = reg_0_2&cdxi2452m;
wire cdxi3195m = reg_0_2&cdxi2453m;
wire cdxi3196m = reg_0_2&cdxi2454m;
wire cdxi3197m = reg_0_1&cdxi2653m;
wire cdxi3198m = reg_0_1&cdxi2654m;
wire cdxi3199m = reg_0_1&cdxi2655m;
wire cdxi3200m = reg_0_1&cdxi2656m;
wire cdxi3201m = reg_0_1&cdxi2657m;
wire cdxi3202m = reg_0_7&cdxi2080m;
wire cdxi3203m = reg_0_6&cdxi3144m;
wire cdxi3204m = reg_0_5&cdxi2152m;
wire cdxi3205m = reg_0_4&cdxi2222m;
wire cdxi3206m = reg_0_2&cdxi2425m;
wire cdxi3207m = reg_0_1&cdxi2627m;
wire cdxi3208m = (cdxi3146m ^ cdxi3147m ^ cdxi3148m ^ cdxi3149m ^ cdxi3150m ^ cdxi3151m ^ cdxi3152m ^ cdxi3153m ^ cdxi3154m ^ cdxi3155m ^ cdxi3156m ^ cdxi3157m ^ cdxi3158m ^ cdxi3159m ^ cdxi3160m ^ cdxi3161m ^ cdxi3162m ^ cdxi3163m ^ cdxi3164m ^ cdxi3165m ^ cdxi3166m ^ cdxi3167m ^ cdxi3168m ^ cdxi3169m ^ cdxi3170m ^ cdxi3171m ^ cdxi3172m ^ cdxi3173m ^ cdxi3174m ^ cdxi3175m ^ cdxi3176m ^ cdxi3177m ^ cdxi3178m ^ cdxi3179m ^ cdxi3180m ^ cdxi3181m ^ cdxi3182m ^ cdxi3183m ^ cdxi3184m ^ cdxi3185m ^ cdxi3186m ^ cdxi3187m ^ cdxi3188m ^ cdxi3189m ^ cdxi3190m ^ cdxi3191m ^ cdxi3192m ^ cdxi3193m ^ cdxi3194m ^ cdxi3195m ^ cdxi3196m ^ cdxi3197m ^ cdxi3198m ^ cdxi3199m ^ cdxi3200m ^ cdxi3201m ^ cdxi3202m ^ cdxi3203m ^ cdxi3204m ^ cdxi3205m ^ cdxi3206m ^ cdxi3207m ^ cdxi3145m);
wire cdxi3209m = reg_0_0&cdxi3208m;
wire cdxi3210m = cdxi1762m&cdxi657m ^ r124m;
wire cdxi3211m = cdxi405m&cdxi1548m;
wire cdxi3212m = cdxi362m&cdxi1232m;
wire cdxi3213m = cdxi362m&cdxi1479m;
wire cdxi3214m = cdxi2256m&cdxi208m;
wire cdxi3215m = cdxi406m&cdxi1549m;
wire cdxi3216m = cdxi362m&cdxi1727m;
wire cdxi3217m = cdxi362m&cdxi1728m;
wire cdxi3218m = cdxi362m&cdxi1729m;
wire cdxi3219m = cdxi362m&cdxi1730m;
wire cdxi3220m = cdxi445m&cdxi1201m;
wire cdxi3221m = cdxi582m&cdxi1273m;
wire cdxi3222m = cdxi1088m&cdxi489m;
wire cdxi3223m = cdxi2323m&r11m;
wire cdxi3224m = cdxi2256m&r12m;
wire cdxi3225m = cdxi446m&cdxi1657m;
wire cdxi3226m = cdxi978m&cdxi623m;
wire cdxi3227m = cdxi406m&cdxi1554m;
wire cdxi3228m = cdxi406m&cdxi1555m;
wire cdxi3229m = cdxi362m&cdxi1731m;
wire cdxi3230m = cdxi362m&cdxi1732m;
wire cdxi3231m = cdxi362m&cdxi1733m;
wire cdxi3232m = cdxi362m&cdxi1734m;
wire cdxi3233m = cdxi362m&cdxi1735m;
wire cdxi3234m = cdxi362m&cdxi1736m;
wire cdxi3235m = cdxi638m&cdxi1135m;
wire cdxi3236m = cdxi466m&cdxi1172m;
wire cdxi3237m = cdxi445m&cdxi1207m;
wire cdxi3238m = cdxi445m&cdxi1208m;
wire cdxi3239m = cdxi1196m&r37m;
wire cdxi3240m = cdxi1160m&r38m;
wire cdxi3241m = cdxi582m&cdxi1280m;
wire cdxi3242m = cdxi1123m&r40m;
wire cdxi3243m = cdxi1088m&r41m;
wire cdxi3244m = cdxi1303m&r42m;
wire cdxi3245m = cdxi1051m&r53m;
wire cdxi3246m = cdxi1161m&r54m;
wire cdxi3247m = cdxi1014m&r55m;
wire cdxi3248m = cdxi1124m&r56m;
wire cdxi3249m = cdxi978m&r57m;
wire cdxi3250m = cdxi1233m&r58m;
wire cdxi3251m = cdxi939m&r59m;
wire cdxi3252m = cdxi901m&r60m;
wire cdxi3253m = cdxi862m&r61m;
wire cdxi3254m = cdxi823m&r62m;
wire cdxi3255m = cdxi657m&r73m;
wire cdxi3256m = cdxi485m&r74m;
wire cdxi3257m = cdxi638m&r75m;
wire cdxi3258m = cdxi562m&r76m;
wire cdxi3259m = cdxi466m&r77m;
wire cdxi3260m = cdxi445m&r78m;
wire cdxi3261m = cdxi425m&r79m;
wire cdxi3262m = cdxi601m&r80m;
wire cdxi3263m = cdxi582m&r81m;
wire cdxi3264m = cdxi405m&r82m;
wire cdxi3265m = cdxi426m&r93m;
wire cdxi3266m = cdxi385m&r94m;
wire cdxi3267m = cdxi446m&r95m;
wire cdxi3268m = cdxi406m&r96m;
wire cdxi3269m = cdxi362m&r97m;
wire cdxi3270m = cdxi207m&r108m;
wire cdxi3271m = cdxi218m&r109m;
wire cdxi3272m = cdxi240m&r110m;
wire cdxi3273m = cdxi196m&r111m;
wire cdxi3274m = cdxi184m&r112m;
wire cdxi3275m = cdxi185m&r118m;
wire cdxi3276m = (cdxi3210m ^ cdxi3214m ^ cdxi3215m ^ cdxi3216m ^ cdxi3217m ^ cdxi3218m ^ cdxi3219m ^ cdxi3220m ^ cdxi3221m ^ cdxi3222m ^ cdxi3223m ^ cdxi3224m ^ cdxi3225m ^ cdxi3226m ^ cdxi3227m ^ cdxi3228m ^ cdxi3229m ^ cdxi3230m ^ cdxi3231m ^ cdxi3232m ^ cdxi3233m ^ cdxi3234m ^ cdxi3235m ^ cdxi3236m ^ cdxi3237m ^ cdxi3238m ^ cdxi3239m ^ cdxi3240m ^ cdxi3241m ^ cdxi3242m ^ cdxi3243m ^ cdxi3244m ^ cdxi3245m ^ cdxi3246m ^ cdxi3247m ^ cdxi3248m ^ cdxi3249m ^ cdxi3250m ^ cdxi3251m ^ cdxi3252m ^ cdxi3253m ^ cdxi3254m ^ cdxi3255m ^ cdxi3256m ^ cdxi3257m ^ cdxi3258m ^ cdxi3259m ^ cdxi3260m ^ cdxi3261m ^ cdxi3262m ^ cdxi3263m ^ cdxi3264m ^ cdxi3265m ^ cdxi3266m ^ cdxi3267m ^ cdxi3268m ^ cdxi3269m ^ cdxi3270m ^ cdxi3271m ^ cdxi3272m ^ cdxi3273m ^ cdxi3274m ^ cdxi3275m);
wire cdxi3277m = a0&cdxi3276m;
wire cdxi3278m = (reg_0_132);
wire cdxi3279m = reg_0_3&cdxi2426m;
wire cdxi3280m = reg_0_1&cdxi2695m;
wire cdxi3281m = reg_0_1&cdxi2696m;
wire cdxi3282m = reg_0_1&cdxi2697m;
wire cdxi3283m = reg_0_1&cdxi2698m;
wire cdxi3284m = reg_0_1&cdxi2699m;
wire cdxi3285m = reg_0_4&reg_0_5&cdxi1219m;
wire cdxi3286m = reg_0_3&cdxi2431m;
wire cdxi3287m = reg_0_3&cdxi2432m;
wire cdxi3288m = reg_0_3&cdxi2433m;
wire cdxi3289m = reg_0_3&cdxi2434m;
wire cdxi3290m = reg_0_1&cdxi2700m;
wire cdxi3291m = reg_0_1&cdxi2701m;
wire cdxi3292m = reg_0_1&cdxi2702m;
wire cdxi3293m = reg_0_1&cdxi2703m;
wire cdxi3294m = reg_0_1&cdxi2704m;
wire cdxi3295m = reg_0_1&cdxi2705m;
wire cdxi3296m = reg_0_1&cdxi2706m;
wire cdxi3297m = reg_0_1&cdxi2707m;
wire cdxi3298m = reg_0_1&cdxi2708m;
wire cdxi3299m = reg_0_1&cdxi2709m;
wire cdxi3300m = reg_0_5&reg_0_6&cdxi1153m;
wire cdxi3301m = reg_0_4&reg_0_6&cdxi1189m;
wire cdxi3302m = reg_0_4&reg_0_5&cdxi1225m;
wire cdxi3303m = reg_0_4&reg_0_5&cdxi1226m;
wire cdxi3304m = reg_0_3&cdxi2441m;
wire cdxi3305m = reg_0_3&cdxi2442m;
wire cdxi3306m = reg_0_3&cdxi2443m;
wire cdxi3307m = reg_0_3&cdxi2444m;
wire cdxi3308m = reg_0_3&cdxi2445m;
wire cdxi3309m = reg_0_3&cdxi2446m;
wire cdxi3310m = reg_0_1&cdxi2710m;
wire cdxi3311m = reg_0_1&cdxi2711m;
wire cdxi3312m = reg_0_1&cdxi2712m;
wire cdxi3313m = reg_0_1&cdxi2713m;
wire cdxi3314m = reg_0_1&cdxi2714m;
wire cdxi3315m = reg_0_1&cdxi2715m;
wire cdxi3316m = reg_0_1&cdxi2716m;
wire cdxi3317m = reg_0_1&cdxi2717m;
wire cdxi3318m = reg_0_1&cdxi2718m;
wire cdxi3319m = reg_0_1&cdxi2719m;
wire cdxi3320m = reg_0_6&cdxi2384m;
wire cdxi3321m = reg_0_5&reg_0_7&cdxi1105m;
wire cdxi3322m = reg_0_5&reg_0_6&cdxi1142m;
wire cdxi3323m = reg_0_4&reg_0_7&cdxi1939m;
wire cdxi3324m = reg_0_4&reg_0_6&cdxi1178m;
wire cdxi3325m = reg_0_4&reg_0_5&cdxi1214m;
wire cdxi3326m = reg_0_3&cdxi2451m;
wire cdxi3327m = reg_0_3&cdxi2452m;
wire cdxi3328m = reg_0_3&cdxi2453m;
wire cdxi3329m = reg_0_3&cdxi2454m;
wire cdxi3330m = reg_0_1&cdxi2720m;
wire cdxi3331m = reg_0_1&cdxi2721m;
wire cdxi3332m = reg_0_1&cdxi2722m;
wire cdxi3333m = reg_0_1&cdxi2723m;
wire cdxi3334m = reg_0_1&cdxi2724m;
wire cdxi3335m = reg_0_7&cdxi2289m;
wire cdxi3336m = reg_0_6&cdxi2358m;
wire cdxi3337m = reg_0_5&cdxi2873m;
wire cdxi3338m = reg_0_4&cdxi3009m;
wire cdxi3339m = reg_0_3&cdxi2425m;
wire cdxi3340m = reg_0_1&cdxi2694m;
wire cdxi3341m = (cdxi3279m ^ cdxi3280m ^ cdxi3281m ^ cdxi3282m ^ cdxi3283m ^ cdxi3284m ^ cdxi3285m ^ cdxi3286m ^ cdxi3287m ^ cdxi3288m ^ cdxi3289m ^ cdxi3290m ^ cdxi3291m ^ cdxi3292m ^ cdxi3293m ^ cdxi3294m ^ cdxi3295m ^ cdxi3296m ^ cdxi3297m ^ cdxi3298m ^ cdxi3299m ^ cdxi3300m ^ cdxi3301m ^ cdxi3302m ^ cdxi3303m ^ cdxi3304m ^ cdxi3305m ^ cdxi3306m ^ cdxi3307m ^ cdxi3308m ^ cdxi3309m ^ cdxi3310m ^ cdxi3311m ^ cdxi3312m ^ cdxi3313m ^ cdxi3314m ^ cdxi3315m ^ cdxi3316m ^ cdxi3317m ^ cdxi3318m ^ cdxi3319m ^ cdxi3320m ^ cdxi3321m ^ cdxi3322m ^ cdxi3323m ^ cdxi3324m ^ cdxi3325m ^ cdxi3326m ^ cdxi3327m ^ cdxi3328m ^ cdxi3329m ^ cdxi3330m ^ cdxi3331m ^ cdxi3332m ^ cdxi3333m ^ cdxi3334m ^ cdxi3335m ^ cdxi3336m ^ cdxi3337m ^ cdxi3338m ^ cdxi3339m ^ cdxi3340m ^ cdxi3278m);
wire cdxi3342m = reg_0_0&cdxi3341m;
wire cdxi3343m = 1&1 ^ cdxi219m ^ cdxi184m ^ cdxi240m ^ cdxi207m;
wire cdxi3344m = cdxi185m&cdxi134m;
wire cdxi3345m = reg_0_1&cdxi137m;
wire cdxi3346m = cdxi219m&cdxi140m;
wire cdxi3347m = reg_0_2&cdxi143m;
wire cdxi3348m = cdxi219m&cdxi146m;
wire cdxi3349m = reg_0_2&cdxi149m;
wire cdxi3350m = cdxi184m&cdxi146m;
wire cdxi3351m = reg_0_3&cdxi149m;
wire cdxi3352m = cdxi196m&cdxi152m;
wire cdxi3353m = reg_0_4&cdxi155m;
wire cdxi3354m = cdxi240m&cdxi168m;
wire cdxi3355m = reg_0_5&cdxi171m;
wire cdxi3356m = cdxi218m&cdxi168m;
wire cdxi3357m = reg_0_6&cdxi171m;
wire cdxi3358m = cdxi363m ^ r7m;
wire cdxi3359m = cdxi219m&r0m;
wire cdxi3360m = cdxi185m&r1m;
wire cdxi3361m = (cdxi3358m ^ cdxi3359m ^ cdxi3360m);
wire cdxi3362m = a0&cdxi3361m;
wire cdxi3363m = reg_0_2&cdxi130m;
wire cdxi3364m = reg_0_1&cdxi136m;
wire cdxi3365m = (cdxi3363m ^ cdxi3364m ^ cdxi372m);
wire cdxi3366m = reg_0_0&cdxi3365m;
wire cdxi3367m = cdxi446m ^ r10m;
wire cdxi3368m = cdxi240m&r0m;
wire cdxi3369m = cdxi185m&r4m;
wire cdxi3370m = (cdxi3367m ^ cdxi3368m ^ cdxi3369m);
wire cdxi3371m = a0&cdxi3370m;
wire cdxi3372m = reg_0_5&cdxi130m;
wire cdxi3373m = reg_0_1&cdxi154m;
wire cdxi3374m = (cdxi3372m ^ cdxi3373m ^ cdxi455m);
wire cdxi3375m = reg_0_0&cdxi3374m;
wire cdxi3376m = cdxi504m ^ r14m;
wire cdxi3377m = cdxi196m&r1m;
wire cdxi3378m = cdxi219m&r3m;
wire cdxi3379m = (cdxi3376m ^ cdxi3377m ^ cdxi3378m);
wire cdxi3380m = a0&cdxi3379m;
wire cdxi3381m = reg_0_4&cdxi136m;
wire cdxi3382m = reg_0_2&cdxi148m;
wire cdxi3383m = (cdxi3381m ^ cdxi3382m ^ cdxi513m);
wire cdxi3384m = reg_0_0&cdxi3383m;
wire cdxi3385m = cdxi524m ^ r15m;
wire cdxi3386m = cdxi240m&r1m;
wire cdxi3387m = cdxi219m&r4m;
wire cdxi3388m = (cdxi3385m ^ cdxi3386m ^ cdxi3387m);
wire cdxi3389m = a0&cdxi3388m;
wire cdxi3390m = reg_0_5&cdxi136m;
wire cdxi3391m = reg_0_2&cdxi154m;
wire cdxi3392m = (cdxi3390m ^ cdxi3391m ^ cdxi533m);
wire cdxi3393m = reg_0_0&cdxi3392m;
wire cdxi3394m = a0&cdxi273m;
wire cdxi3395m = reg_0_0&cdxi278m;
wire cdxi3396m = a0&cdxi283m;
wire cdxi3397m = reg_0_0&cdxi288m;
wire cdxi3398m = a0&cdxi313m;
wire cdxi3399m = reg_0_0&cdxi318m;
wire cdxi3400m = a0&cdxi303m;
wire cdxi3401m = reg_0_0&cdxi308m;
wire cdxi3402m = a0&cdxi327m;
wire cdxi3403m = reg_0_0&cdxi332m;
wire cdxi3404m = a0&cdxi339m;
wire cdxi3405m = reg_0_0&cdxi344m;
wire cdxi3406m = cdxi185m&cdxi3379m;
wire cdxi3407m = reg_0_1&cdxi3383m;
wire cdxi3408m = cdxi185m&cdxi3388m;
wire cdxi3409m = reg_0_1&cdxi3392m;
wire cdxi3410m = cdxi185m&cdxi327m;
wire cdxi3411m = reg_0_1&cdxi332m;
wire cdxi3412m = cdxi219m&cdxi283m;
wire cdxi3413m = reg_0_2&cdxi288m;
wire cdxi3414m = cdxi219m&cdxi293m;
wire cdxi3415m = reg_0_2&cdxi298m;
wire cdxi3416m = cdxi219m&cdxi243m;
wire cdxi3417m = reg_0_2&cdxi248m;
wire cdxi3418m = cdxi219m&cdxi263m;
wire cdxi3419m = reg_0_2&cdxi268m;
wire cdxi3420m = cdxi240m&cdxi339m;
wire cdxi3421m = reg_0_5&cdxi344m;
wire cdxi3422m = cdxi824m ^ r29m;
wire cdxi3423m = cdxi219m&cdxi197m;
wire cdxi3424m = cdxi406m&r1m;
wire cdxi3425m = cdxi363m&r3m;
wire cdxi3426m = cdxi196m&r7m;
wire cdxi3427m = cdxi219m&r9m;
wire cdxi3428m = cdxi185m&r14m;
wire cdxi3429m = (cdxi3422m ^ cdxi3423m ^ cdxi3424m ^ cdxi3425m ^ cdxi3426m ^ cdxi3427m ^ cdxi3428m);
wire cdxi3430m = a0&cdxi3429m;
wire cdxi3431m = reg_0_2&cdxi202m;
wire cdxi3432m = reg_0_1&cdxi3381m;
wire cdxi3433m = reg_0_1&cdxi3382m;
wire cdxi3434m = reg_0_4&cdxi372m;
wire cdxi3435m = reg_0_2&cdxi201m;
wire cdxi3436m = reg_0_1&cdxi513m;
wire cdxi3437m = (cdxi3431m ^ cdxi3432m ^ cdxi3433m ^ cdxi3434m ^ cdxi3435m ^ cdxi3436m ^ cdxi842m);
wire cdxi3438m = reg_0_0&cdxi3437m;
wire cdxi3439m = cdxi940m ^ r32m;
wire cdxi3440m = cdxi219m&cdxi208m;
wire cdxi3441m = cdxi185m&cdxi271m;
wire cdxi3442m = cdxi185m&cdxi272m;
wire cdxi3443m = cdxi207m&r7m;
wire cdxi3444m = cdxi219m&r12m;
wire cdxi3445m = cdxi185m&r17m;
wire cdxi3446m = (cdxi3439m ^ cdxi3440m ^ cdxi3441m ^ cdxi3442m ^ cdxi3443m ^ cdxi3444m ^ cdxi3445m);
wire cdxi3447m = a0&cdxi3446m;
wire cdxi3448m = reg_0_2&cdxi213m;
wire cdxi3449m = reg_0_1&cdxi276m;
wire cdxi3450m = reg_0_1&cdxi277m;
wire cdxi3451m = reg_0_7&cdxi372m;
wire cdxi3452m = reg_0_2&cdxi212m;
wire cdxi3453m = reg_0_1&cdxi275m;
wire cdxi3454m = (cdxi3448m ^ cdxi3449m ^ cdxi3450m ^ cdxi3451m ^ cdxi3452m ^ cdxi3453m ^ cdxi957m);
wire cdxi3455m = reg_0_0&cdxi3454m;
wire cdxi3456m = cdxi862m ^ r34m;
wire cdxi3457m = cdxi582m&r0m;
wire cdxi3458m = cdxi185m&cdxi311m;
wire cdxi3459m = cdxi185m&cdxi312m;
wire cdxi3460m = cdxi240m&r8m;
wire cdxi3461m = cdxi184m&r10m;
wire cdxi3462m = cdxi185m&r19m;
wire cdxi3463m = (cdxi3456m ^ cdxi3457m ^ cdxi3458m ^ cdxi3459m ^ cdxi3460m ^ cdxi3461m ^ cdxi3462m);
wire cdxi3464m = a0&cdxi3463m;
wire cdxi3465m = reg_0_3&cdxi3372m;
wire cdxi3466m = reg_0_1&cdxi316m;
wire cdxi3467m = reg_0_1&cdxi317m;
wire cdxi3468m = reg_0_5&cdxi190m;
wire cdxi3469m = reg_0_3&cdxi455m;
wire cdxi3470m = reg_0_1&cdxi315m;
wire cdxi3471m = (cdxi3465m ^ cdxi3466m ^ cdxi3467m ^ cdxi3468m ^ cdxi3469m ^ cdxi3470m ^ cdxi881m);
wire cdxi3472m = reg_0_0&cdxi3471m;
wire cdxi3473m = cdxi901m ^ r35m;
wire cdxi3474m = cdxi601m&r0m;
wire cdxi3475m = cdxi185m&cdxi291m;
wire cdxi3476m = cdxi185m&cdxi292m;
wire cdxi3477m = cdxi218m&r8m;
wire cdxi3478m = cdxi184m&r11m;
wire cdxi3479m = cdxi185m&r20m;
wire cdxi3480m = (cdxi3473m ^ cdxi3474m ^ cdxi3475m ^ cdxi3476m ^ cdxi3477m ^ cdxi3478m ^ cdxi3479m);
wire cdxi3481m = a0&cdxi3480m;
wire cdxi3482m = reg_0_3&reg_0_6&cdxi130m;
wire cdxi3483m = reg_0_1&cdxi296m;
wire cdxi3484m = reg_0_1&cdxi297m;
wire cdxi3485m = reg_0_6&cdxi190m;
wire cdxi3486m = reg_0_3&cdxi394m;
wire cdxi3487m = reg_0_1&cdxi295m;
wire cdxi3488m = (cdxi3482m ^ cdxi3483m ^ cdxi3484m ^ cdxi3485m ^ cdxi3486m ^ cdxi3487m ^ cdxi919m);
wire cdxi3489m = reg_0_0&cdxi3488m;
wire cdxi3490m = a0&cdxi700m;
wire cdxi3491m = reg_0_0&cdxi709m;
wire cdxi3492m = cdxi938m ^ r46m;
wire cdxi3493m = cdxi184m&cdxi271m;
wire cdxi3494m = cdxi219m&cdxi230m;
wire cdxi3495m = cdxi219m&cdxi231m;
wire cdxi3496m = cdxi207m&r13m;
wire cdxi3497m = cdxi184m&r17m;
wire cdxi3498m = cdxi219m&r21m;
wire cdxi3499m = (cdxi3492m ^ cdxi3493m ^ cdxi3494m ^ cdxi3495m ^ cdxi3496m ^ cdxi3497m ^ cdxi3498m);
wire cdxi3500m = a0&cdxi3499m;
wire cdxi3501m = reg_0_3&cdxi276m;
wire cdxi3502m = reg_0_2&cdxi235m;
wire cdxi3503m = reg_0_2&cdxi236m;
wire cdxi3504m = reg_0_7&cdxi373m;
wire cdxi3505m = reg_0_3&cdxi275m;
wire cdxi3506m = reg_0_2&cdxi234m;
wire cdxi3507m = (cdxi3501m ^ cdxi3502m ^ cdxi3503m ^ cdxi3504m ^ cdxi3505m ^ cdxi3506m ^ cdxi958m);
wire cdxi3508m = reg_0_0&cdxi3507m;
wire cdxi3509m = cdxi1050m ^ r52m;
wire cdxi3510m = cdxi218m&cdxi271m;
wire cdxi3511m = cdxi219m&cdxi337m;
wire cdxi3512m = cdxi219m&cdxi338m;
wire cdxi3513m = cdxi207m&r16m;
wire cdxi3514m = cdxi218m&r17m;
wire cdxi3515m = cdxi219m&r27m;
wire cdxi3516m = (cdxi3509m ^ cdxi3510m ^ cdxi3511m ^ cdxi3512m ^ cdxi3513m ^ cdxi3514m ^ cdxi3515m);
wire cdxi3517m = a0&cdxi3516m;
wire cdxi3518m = reg_0_6&cdxi276m;
wire cdxi3519m = reg_0_2&cdxi342m;
wire cdxi3520m = reg_0_2&cdxi343m;
wire cdxi3521m = reg_0_7&cdxi224m;
wire cdxi3522m = reg_0_6&cdxi275m;
wire cdxi3523m = reg_0_2&cdxi341m;
wire cdxi3524m = (cdxi3518m ^ cdxi3519m ^ cdxi3520m ^ cdxi3521m ^ cdxi3522m ^ cdxi3523m ^ cdxi1069m);
wire cdxi3525m = reg_0_0&cdxi3524m;
wire cdxi3526m = a0&cdxi784m;
wire cdxi3527m = reg_0_0&cdxi793m;
wire cdxi3528m = cdxi1374m ^ r56m;
wire cdxi3529m = cdxi240m&cdxi291m;
wire cdxi3530m = cdxi184m&cdxi251m;
wire cdxi3531m = cdxi184m&cdxi252m;
wire cdxi3532m = cdxi218m&r19m;
wire cdxi3533m = cdxi240m&r20m;
wire cdxi3534m = cdxi184m&r25m;
wire cdxi3535m = (cdxi3528m ^ cdxi3529m ^ cdxi3530m ^ cdxi3531m ^ cdxi3532m ^ cdxi3533m ^ cdxi3534m);
wire cdxi3536m = a0&cdxi3535m;
wire cdxi3537m = reg_0_5&cdxi296m;
wire cdxi3538m = reg_0_3&cdxi256m;
wire cdxi3539m = reg_0_3&cdxi257m;
wire cdxi3540m = reg_0_6&cdxi315m;
wire cdxi3541m = reg_0_5&cdxi295m;
wire cdxi3542m = reg_0_3&cdxi255m;
wire cdxi3543m = (cdxi3537m ^ cdxi3538m ^ cdxi3539m ^ cdxi3540m ^ cdxi3541m ^ cdxi3542m ^ cdxi1391m);
wire cdxi3544m = reg_0_0&cdxi3543m;
wire cdxi3545m = a0&cdxi808m;
wire cdxi3546m = reg_0_0&cdxi817m;
wire cdxi3547m = cdxi185m&cdxi511m;
wire cdxi3548m = reg_0_1&cdxi521m;
wire cdxi3549m = cdxi185m&cdxi3499m;
wire cdxi3550m = reg_0_1&cdxi3507m;
wire cdxi3551m = cdxi185m&cdxi3516m;
wire cdxi3552m = reg_0_1&cdxi3524m;
wire cdxi3553m = cdxi185m&cdxi784m;
wire cdxi3554m = reg_0_1&cdxi793m;
wire cdxi3555m = cdxi185m&cdxi3535m;
wire cdxi3556m = reg_0_1&cdxi3543m;
wire cdxi3557m = cdxi185m&cdxi664m;
wire cdxi3558m = reg_0_1&cdxi673m;
wire cdxi3559m = cdxi219m&cdxi608m;
wire cdxi3560m = reg_0_2&cdxi617m;
wire cdxi3561m = cdxi1196m ^ r58m;
wire cdxi3562m = cdxi218m&cdxi230m;
wire cdxi3563m = cdxi184m&cdxi337m;
wire cdxi3564m = cdxi184m&cdxi338m;
wire cdxi3565m = cdxi207m&r20m;
wire cdxi3566m = cdxi218m&r21m;
wire cdxi3567m = cdxi184m&r27m;
wire cdxi3568m = (cdxi3561m ^ cdxi3562m ^ cdxi3563m ^ cdxi3564m ^ cdxi3565m ^ cdxi3566m ^ cdxi3567m);
wire cdxi3569m = cdxi219m&cdxi3568m;
wire cdxi3570m = reg_0_6&cdxi235m;
wire cdxi3571m = reg_0_3&cdxi342m;
wire cdxi3572m = reg_0_3&cdxi343m;
wire cdxi3573m = reg_0_7&cdxi295m;
wire cdxi3574m = reg_0_6&cdxi234m;
wire cdxi3575m = reg_0_3&cdxi341m;
wire cdxi3576m = (cdxi3570m ^ cdxi3571m ^ cdxi3572m ^ cdxi3573m ^ cdxi3574m ^ cdxi3575m ^ cdxi1213m);
wire cdxi3577m = reg_0_2&cdxi3576m;
wire cdxi3578m = cdxi219m&cdxi808m;
wire cdxi3579m = reg_0_2&cdxi817m;
wire cdxi3580m = cdxi184m&cdxi664m;
wire cdxi3581m = reg_0_3&cdxi673m;
wire cdxi3582m = cdxi196m&cdxi664m;
wire cdxi3583m = reg_0_4&cdxi673m;
wire cdxi3584m = cdxi2117m ^ r69m;
wire cdxi3585m = cdxi504m&cdxi208m;
wire cdxi3586m = cdxi406m&cdxi271m;
wire cdxi3587m = cdxi363m&cdxi325m;
wire cdxi3588m = cdxi363m&cdxi326m;
wire cdxi3589m = cdxi562m&r7m;
wire cdxi3590m = cdxi563m&r9m;
wire cdxi3591m = cdxi504m&r12m;
wire cdxi3592m = cdxi426m&r14m;
wire cdxi3593m = cdxi406m&r17m;
wire cdxi3594m = cdxi363m&r24m;
wire cdxi3595m = cdxi207m&r29m;
wire cdxi3596m = cdxi196m&r32m;
wire cdxi3597m = cdxi219m&r39m;
wire cdxi3598m = cdxi185m&r49m;
wire cdxi3599m = (cdxi3584m ^ cdxi3585m ^ cdxi3586m ^ cdxi3587m ^ cdxi3588m ^ cdxi3589m ^ cdxi3590m ^ cdxi3591m ^ cdxi3592m ^ cdxi3593m ^ cdxi3594m ^ cdxi3595m ^ cdxi3596m ^ cdxi3597m ^ cdxi3598m);
wire cdxi3600m = a0&cdxi3599m;
wire cdxi3601m = reg_0_2&reg_0_4&cdxi213m;
wire cdxi3602m = reg_0_1&cdxi573m;
wire cdxi3603m = reg_0_1&cdxi574m;
wire cdxi3604m = reg_0_1&cdxi575m;
wire cdxi3605m = reg_0_4&cdxi3451m;
wire cdxi3606m = reg_0_2&reg_0_7&cdxi201m;
wire cdxi3607m = reg_0_2&reg_0_4&cdxi212m;
wire cdxi3608m = reg_0_1&cdxi576m;
wire cdxi3609m = reg_0_1&cdxi577m;
wire cdxi3610m = reg_0_1&cdxi578m;
wire cdxi3611m = reg_0_7&cdxi842m;
wire cdxi3612m = reg_0_4&cdxi957m;
wire cdxi3613m = reg_0_2&cdxi1141m;
wire cdxi3614m = reg_0_1&cdxi572m;
wire cdxi3615m = (cdxi3601m ^ cdxi3602m ^ cdxi3603m ^ cdxi3604m ^ cdxi3605m ^ cdxi3606m ^ cdxi3607m ^ cdxi3608m ^ cdxi3609m ^ cdxi3610m ^ cdxi3611m ^ cdxi3612m ^ cdxi3613m ^ cdxi3614m ^ cdxi2150m);
wire cdxi3616m = reg_0_0&cdxi3615m;
wire cdxi3617m = cdxi2187m ^ r82m;
wire cdxi3618m = cdxi638m&cdxi208m;
wire cdxi3619m = cdxi385m&cdxi261m;
wire cdxi3620m = cdxi446m&cdxi337m;
wire cdxi3621m = cdxi446m&cdxi338m;
wire cdxi3622m = cdxi218m&cdxi489m;
wire cdxi3623m = cdxi485m&r11m;
wire cdxi3624m = cdxi638m&r12m;
wire cdxi3625m = cdxi426m&r25m;
wire cdxi3626m = cdxi385m&r26m;
wire cdxi3627m = cdxi446m&r27m;
wire cdxi3628m = cdxi207m&r40m;
wire cdxi3629m = cdxi218m&r41m;
wire cdxi3630m = cdxi240m&r42m;
wire cdxi3631m = cdxi185m&r62m;
wire cdxi3632m = (cdxi3617m ^ cdxi3618m ^ cdxi3619m ^ cdxi3620m ^ cdxi3621m ^ cdxi3622m ^ cdxi3623m ^ cdxi3624m ^ cdxi3625m ^ cdxi3626m ^ cdxi3627m ^ cdxi3628m ^ cdxi3629m ^ cdxi3630m ^ cdxi3631m);
wire cdxi3633m = a0&cdxi3632m;
wire cdxi3634m = reg_0_5&reg_0_6&cdxi213m;
wire cdxi3635m = reg_0_1&cdxi667m;
wire cdxi3636m = reg_0_1&cdxi668m;
wire cdxi3637m = reg_0_1&cdxi669m;
wire cdxi3638m = reg_0_6&cdxi498m;
wire cdxi3639m = reg_0_5&reg_0_7&cdxi394m;
wire cdxi3640m = reg_0_5&reg_0_6&cdxi212m;
wire cdxi3641m = reg_0_1&cdxi670m;
wire cdxi3642m = reg_0_1&cdxi671m;
wire cdxi3643m = reg_0_1&cdxi672m;
wire cdxi3644m = reg_0_7&cdxi1031m;
wire cdxi3645m = reg_0_6&cdxi494m;
wire cdxi3646m = reg_0_5&cdxi1068m;
wire cdxi3647m = reg_0_1&cdxi666m;
wire cdxi3648m = (cdxi3634m ^ cdxi3635m ^ cdxi3636m ^ cdxi3637m ^ cdxi3638m ^ cdxi3639m ^ cdxi3640m ^ cdxi3641m ^ cdxi3642m ^ cdxi3643m ^ cdxi3644m ^ cdxi3645m ^ cdxi3646m ^ cdxi3647m ^ cdxi2220m);
wire cdxi3649m = reg_0_0&cdxi3648m;
wire cdxi3650m = cdxi2114m ^ r91m;
wire cdxi3651m = cdxi466m&cdxi271m;
wire cdxi3652m = cdxi384m&cdxi325m;
wire cdxi3653m = cdxi504m&cdxi337m;
wire cdxi3654m = cdxi504m&cdxi338m;
wire cdxi3655m = cdxi218m&cdxi567m;
wire cdxi3656m = cdxi562m&r16m;
wire cdxi3657m = cdxi466m&r17m;
wire cdxi3658m = cdxi563m&r23m;
wire cdxi3659m = cdxi384m&r24m;
wire cdxi3660m = cdxi504m&r27m;
wire cdxi3661m = cdxi207m&r48m;
wire cdxi3662m = cdxi218m&r49m;
wire cdxi3663m = cdxi196m&r52m;
wire cdxi3664m = cdxi219m&r61m;
wire cdxi3665m = (cdxi3650m ^ cdxi3651m ^ cdxi3652m ^ cdxi3653m ^ cdxi3654m ^ cdxi3655m ^ cdxi3656m ^ cdxi3657m ^ cdxi3658m ^ cdxi3659m ^ cdxi3660m ^ cdxi3661m ^ cdxi3662m ^ cdxi3663m ^ cdxi3664m);
wire cdxi3666m = a0&cdxi3665m;
wire cdxi3667m = reg_0_4&cdxi3518m;
wire cdxi3668m = reg_0_2&cdxi767m;
wire cdxi3669m = reg_0_2&cdxi768m;
wire cdxi3670m = reg_0_2&cdxi769m;
wire cdxi3671m = reg_0_6&cdxi576m;
wire cdxi3672m = reg_0_4&cdxi3521m;
wire cdxi3673m = reg_0_4&cdxi3522m;
wire cdxi3674m = reg_0_2&cdxi770m;
wire cdxi3675m = reg_0_2&cdxi771m;
wire cdxi3676m = reg_0_2&cdxi772m;
wire cdxi3677m = reg_0_7&cdxi552m;
wire cdxi3678m = reg_0_6&cdxi572m;
wire cdxi3679m = reg_0_4&cdxi1069m;
wire cdxi3680m = reg_0_2&cdxi766m;
wire cdxi3681m = (cdxi3667m ^ cdxi3668m ^ cdxi3669m ^ cdxi3670m ^ cdxi3671m ^ cdxi3672m ^ cdxi3673m ^ cdxi3674m ^ cdxi3675m ^ cdxi3676m ^ cdxi3677m ^ cdxi3678m ^ cdxi3679m ^ cdxi3680m ^ cdxi2151m);
wire cdxi3682m = reg_0_0&cdxi3681m;
wire cdxi3683m = cdxi2186m ^ r92m;
wire cdxi3684m = cdxi638m&cdxi271m;
wire cdxi3685m = cdxi384m&cdxi261m;
wire cdxi3686m = cdxi524m&cdxi337m;
wire cdxi3687m = cdxi524m&cdxi338m;
wire cdxi3688m = cdxi657m&r15m;
wire cdxi3689m = cdxi485m&r16m;
wire cdxi3690m = cdxi638m&r17m;
wire cdxi3691m = cdxi563m&r25m;
wire cdxi3692m = cdxi384m&r26m;
wire cdxi3693m = cdxi524m&r27m;
wire cdxi3694m = cdxi207m&r50m;
wire cdxi3695m = cdxi218m&r51m;
wire cdxi3696m = cdxi240m&r52m;
wire cdxi3697m = cdxi219m&r62m;
wire cdxi3698m = (cdxi3683m ^ cdxi3684m ^ cdxi3685m ^ cdxi3686m ^ cdxi3687m ^ cdxi3688m ^ cdxi3689m ^ cdxi3690m ^ cdxi3691m ^ cdxi3692m ^ cdxi3693m ^ cdxi3694m ^ cdxi3695m ^ cdxi3696m ^ cdxi3697m);
wire cdxi3699m = a0&cdxi3698m;
wire cdxi3700m = reg_0_5&cdxi3518m;
wire cdxi3701m = reg_0_2&cdxi667m;
wire cdxi3702m = reg_0_2&cdxi668m;
wire cdxi3703m = reg_0_2&cdxi669m;
wire cdxi3704m = reg_0_6&cdxi746m;
wire cdxi3705m = reg_0_5&cdxi3521m;
wire cdxi3706m = reg_0_5&cdxi3522m;
wire cdxi3707m = reg_0_2&cdxi670m;
wire cdxi3708m = reg_0_2&cdxi671m;
wire cdxi3709m = reg_0_2&cdxi672m;
wire cdxi3710m = reg_0_7&cdxi724m;
wire cdxi3711m = reg_0_6&cdxi742m;
wire cdxi3712m = reg_0_5&cdxi1069m;
wire cdxi3713m = reg_0_2&cdxi666m;
wire cdxi3714m = (cdxi3700m ^ cdxi3701m ^ cdxi3702m ^ cdxi3703m ^ cdxi3704m ^ cdxi3705m ^ cdxi3706m ^ cdxi3707m ^ cdxi3708m ^ cdxi3709m ^ cdxi3710m ^ cdxi3711m ^ cdxi3712m ^ cdxi3713m ^ cdxi2221m);
wire cdxi3715m = reg_0_0&cdxi3714m;
wire cdxi3716m = a0&cdxi1667m;
wire cdxi3717m = reg_0_0&cdxi1684m;
wire cdxi3718m = a0&cdxi1741m;
wire cdxi3719m = reg_0_0&cdxi1758m;
wire cdxi3720m = cdxi185m&cdxi1319m;
wire cdxi3721m = reg_0_1&cdxi1336m;
wire cdxi3722m = cdxi185m&cdxi1389m;
wire cdxi3723m = reg_0_1&cdxi1407m;
wire cdxi3724m = cdxi185m&cdxi1425m;
wire cdxi3725m = reg_0_1&cdxi1442m;
wire cdxi3726m = cdxi185m&cdxi3698m;
wire cdxi3727m = reg_0_1&cdxi3714m;
wire cdxi3728m = cdxi185m&cdxi1563m;
wire cdxi3729m = reg_0_1&cdxi1580m;
wire cdxi3730m = cdxi185m&cdxi1741m;
wire cdxi3731m = reg_0_1&cdxi1758m;
wire cdxi3732m = cdxi219m&cdxi1741m;
wire cdxi3733m = reg_0_2&cdxi1758m;
wire cdxi3734m = cdxi2803m ^ r103m;
wire cdxi3735m = cdxi900m&cdxi208m;
wire cdxi3736m = cdxi901m&cdxi271m;
wire cdxi3737m = cdxi902m&cdxi230m;
wire cdxi3738m = cdxi825m&cdxi337m;
wire cdxi3739m = cdxi825m&cdxi338m;
wire cdxi3740m = cdxi1196m&r7m;
wire cdxi3741m = cdxi384m&cdxi430m;
wire cdxi3742m = cdxi938m&r11m;
wire cdxi3743m = cdxi900m&r12m;
wire cdxi3744m = cdxi1051m&r13m;
wire cdxi3745m = cdxi939m&r16m;
wire cdxi3746m = cdxi901m&r17m;
wire cdxi3747m = cdxi940m&r20m;
wire cdxi3748m = cdxi902m&r21m;
wire cdxi3749m = cdxi825m&r27m;
wire cdxi3750m = cdxi657m&r28m;
wire cdxi3751m = cdxi425m&r31m;
wire cdxi3752m = cdxi601m&r32m;
wire cdxi3753m = cdxi563m&r35m;
wire cdxi3754m = cdxi384m&r36m;
wire cdxi3755m = cdxi361m&r42m;
wire cdxi3756m = cdxi426m&r45m;
wire cdxi3757m = cdxi385m&r46m;
wire cdxi3758m = cdxi362m&r52m;
wire cdxi3759m = cdxi363m&r58m;
wire cdxi3760m = cdxi207m&r65m;
wire cdxi3761m = cdxi218m&r66m;
wire cdxi3762m = cdxi184m&r72m;
wire cdxi3763m = cdxi219m&r78m;
wire cdxi3764m = cdxi185m&r88m;
wire cdxi3765m = (cdxi3734m ^ cdxi3735m ^ cdxi3736m ^ cdxi3737m ^ cdxi3738m ^ cdxi3739m ^ cdxi3740m ^ cdxi3741m ^ cdxi3742m ^ cdxi3743m ^ cdxi3744m ^ cdxi3745m ^ cdxi3746m ^ cdxi3747m ^ cdxi3748m ^ cdxi3749m ^ cdxi3750m ^ cdxi3751m ^ cdxi3752m ^ cdxi3753m ^ cdxi3754m ^ cdxi3755m ^ cdxi3756m ^ cdxi3757m ^ cdxi3758m ^ cdxi3759m ^ cdxi3760m ^ cdxi3761m ^ cdxi3762m ^ cdxi3763m ^ cdxi3764m);
wire cdxi3766m = a0&cdxi3765m;
wire cdxi3767m = reg_0_2&cdxi1215m;
wire cdxi3768m = reg_0_1&cdxi1462m;
wire cdxi3769m = reg_0_1&cdxi1463m;
wire cdxi3770m = reg_0_1&cdxi1464m;
wire cdxi3771m = reg_0_1&cdxi1465m;
wire cdxi3772m = reg_0_3&cdxi1075m;
wire cdxi3773m = reg_0_2&cdxi1219m;
wire cdxi3774m = reg_0_2&cdxi1220m;
wire cdxi3775m = reg_0_2&cdxi1221m;
wire cdxi3776m = reg_0_1&cdxi1466m;
wire cdxi3777m = reg_0_1&cdxi1467m;
wire cdxi3778m = reg_0_1&cdxi1468m;
wire cdxi3779m = reg_0_1&cdxi1469m;
wire cdxi3780m = reg_0_1&cdxi1470m;
wire cdxi3781m = reg_0_1&cdxi1471m;
wire cdxi3782m = reg_0_6&cdxi970m;
wire cdxi3783m = reg_0_3&cdxi1081m;
wire cdxi3784m = reg_0_3&cdxi1082m;
wire cdxi3785m = reg_0_2&cdxi1225m;
wire cdxi3786m = reg_0_2&cdxi1226m;
wire cdxi3787m = reg_0_2&cdxi1227m;
wire cdxi3788m = reg_0_1&cdxi1472m;
wire cdxi3789m = reg_0_1&cdxi1473m;
wire cdxi3790m = reg_0_1&cdxi1474m;
wire cdxi3791m = reg_0_1&cdxi1475m;
wire cdxi3792m = reg_0_7&cdxi920m;
wire cdxi3793m = reg_0_6&cdxi959m;
wire cdxi3794m = reg_0_3&cdxi1070m;
wire cdxi3795m = reg_0_2&cdxi1214m;
wire cdxi3796m = reg_0_1&cdxi1461m;
wire cdxi3797m = (cdxi3767m ^ cdxi3768m ^ cdxi3769m ^ cdxi3770m ^ cdxi3771m ^ cdxi3772m ^ cdxi3773m ^ cdxi3774m ^ cdxi3775m ^ cdxi3776m ^ cdxi3777m ^ cdxi3778m ^ cdxi3779m ^ cdxi3780m ^ cdxi3781m ^ cdxi3782m ^ cdxi3783m ^ cdxi3784m ^ cdxi3785m ^ cdxi3786m ^ cdxi3787m ^ cdxi3788m ^ cdxi3789m ^ cdxi3790m ^ cdxi3791m ^ cdxi3792m ^ cdxi3793m ^ cdxi3794m ^ cdxi3795m ^ cdxi3796m ^ cdxi2872m);
wire cdxi3798m = reg_0_0&cdxi3797m;
wire cdxi3799m = cdxi361m&cdxi1479m ^ r113m;
wire cdxi3800m = cdxi405m&cdxi716m;
wire cdxi3801m = cdxi1304m&cdxi291m;
wire cdxi3802m = cdxi361m&cdxi639m;
wire cdxi3803m = cdxi361m&cdxi640m;
wire cdxi3804m = cdxi361m&cdxi641m;
wire cdxi3805m = cdxi445m&cdxi697m;
wire cdxi3806m = cdxi582m&cdxi547m;
wire cdxi3807m = cdxi405m&cdxi719m;
wire cdxi3808m = cdxi405m&cdxi720m;
wire cdxi3809m = cdxi524m&cdxi605m;
wire cdxi3810m = cdxi977m&r19m;
wire cdxi3811m = cdxi1304m&r20m;
wire cdxi3812m = cdxi361m&cdxi642m;
wire cdxi3813m = cdxi361m&cdxi643m;
wire cdxi3814m = cdxi361m&cdxi644m;
wire cdxi3815m = cdxi638m&r43m;
wire cdxi3816m = cdxi466m&r44m;
wire cdxi3817m = cdxi445m&r45m;
wire cdxi3818m = cdxi601m&r47m;
wire cdxi3819m = cdxi582m&r48m;
wire cdxi3820m = cdxi405m&r50m;
wire cdxi3821m = cdxi384m&r53m;
wire cdxi3822m = cdxi524m&r54m;
wire cdxi3823m = cdxi504m&r56m;
wire cdxi3824m = cdxi361m&r59m;
wire cdxi3825m = cdxi218m&r83m;
wire cdxi3826m = cdxi240m&r84m;
wire cdxi3827m = cdxi196m&r86m;
wire cdxi3828m = cdxi184m&r89m;
wire cdxi3829m = cdxi219m&r93m;
wire cdxi3830m = (cdxi3799m ^ cdxi3800m ^ cdxi3801m ^ cdxi3802m ^ cdxi3803m ^ cdxi3804m ^ cdxi3805m ^ cdxi3806m ^ cdxi3807m ^ cdxi3808m ^ cdxi3809m ^ cdxi3810m ^ cdxi3811m ^ cdxi3812m ^ cdxi3813m ^ cdxi3814m ^ cdxi3815m ^ cdxi3816m ^ cdxi3817m ^ cdxi3818m ^ cdxi3819m ^ cdxi3820m ^ cdxi3821m ^ cdxi3822m ^ cdxi3823m ^ cdxi3824m ^ cdxi3825m ^ cdxi3826m ^ cdxi3827m ^ cdxi3828m ^ cdxi3829m);
wire cdxi3831m = a0&cdxi3830m;
wire cdxi3832m = (reg_0_121);
wire cdxi3833m = reg_0_3&cdxi1497m;
wire cdxi3834m = reg_0_2&cdxi1704m;
wire cdxi3835m = reg_0_2&cdxi1705m;
wire cdxi3836m = reg_0_2&cdxi1706m;
wire cdxi3837m = reg_0_2&cdxi1707m;
wire cdxi3838m = reg_0_4&cdxi1397m;
wire cdxi3839m = reg_0_3&cdxi1501m;
wire cdxi3840m = reg_0_3&cdxi1502m;
wire cdxi3841m = reg_0_3&cdxi1503m;
wire cdxi3842m = reg_0_2&cdxi1708m;
wire cdxi3843m = reg_0_2&cdxi1709m;
wire cdxi3844m = reg_0_2&cdxi1710m;
wire cdxi3845m = reg_0_2&cdxi1711m;
wire cdxi3846m = reg_0_2&cdxi1712m;
wire cdxi3847m = reg_0_2&cdxi1713m;
wire cdxi3848m = reg_0_5&cdxi1610m;
wire cdxi3849m = reg_0_4&cdxi1403m;
wire cdxi3850m = reg_0_4&cdxi1404m;
wire cdxi3851m = reg_0_3&cdxi1507m;
wire cdxi3852m = reg_0_3&cdxi1508m;
wire cdxi3853m = reg_0_3&cdxi1509m;
wire cdxi3854m = reg_0_2&cdxi1714m;
wire cdxi3855m = reg_0_2&cdxi1715m;
wire cdxi3856m = reg_0_2&cdxi1716m;
wire cdxi3857m = reg_0_2&cdxi1717m;
wire cdxi3858m = reg_0_6&cdxi1321m;
wire cdxi3859m = reg_0_5&cdxi1599m;
wire cdxi3860m = reg_0_4&cdxi1392m;
wire cdxi3861m = reg_0_3&cdxi1496m;
wire cdxi3862m = reg_0_2&cdxi1703m;
wire cdxi3863m = (cdxi3833m ^ cdxi3834m ^ cdxi3835m ^ cdxi3836m ^ cdxi3837m ^ cdxi3838m ^ cdxi3839m ^ cdxi3840m ^ cdxi3841m ^ cdxi3842m ^ cdxi3843m ^ cdxi3844m ^ cdxi3845m ^ cdxi3846m ^ cdxi3847m ^ cdxi3848m ^ cdxi3849m ^ cdxi3850m ^ cdxi3851m ^ cdxi3852m ^ cdxi3853m ^ cdxi3854m ^ cdxi3855m ^ cdxi3856m ^ cdxi3857m ^ cdxi3858m ^ cdxi3859m ^ cdxi3860m ^ cdxi3861m ^ cdxi3862m ^ cdxi3832m);
wire cdxi3864m = reg_0_0&cdxi3863m;
wire cdxi3865m = cdxi825m&cdxi1479m ^ r119m;
wire cdxi3866m = cdxi361m&cdxi1479m;
wire cdxi3867m = cdxi825m&cdxi445m;
wire cdxi3868m = cdxi3866m&r0m;
wire cdxi3869m = cdxi362m&cdxi1480m;
wire cdxi3870m = cdxi363m&cdxi1687m;
wire cdxi3871m = cdxi825m&cdxi639m;
wire cdxi3872m = cdxi825m&cdxi640m;
wire cdxi3873m = cdxi825m&cdxi641m;
wire cdxi3874m = cdxi405m&cdxi1019m;
wire cdxi3875m = cdxi2045m&r8m;
wire cdxi3876m = cdxi861m&cdxi470m;
wire cdxi3877m = cdxi1834m&r10m;
wire cdxi3878m = cdxi1761m&r11m;
wire cdxi3879m = cdxi406m&cdxi1379m;
wire cdxi3880m = cdxi862m&cdxi547m;
wire cdxi3881m = cdxi362m&cdxi1485m;
wire cdxi3882m = cdxi362m&cdxi1486m;
wire cdxi3883m = cdxi863m&cdxi605m;
wire cdxi3884m = cdxi363m&cdxi1692m;
wire cdxi3885m = cdxi363m&cdxi1693m;
wire cdxi3886m = cdxi825m&cdxi642m;
wire cdxi3887m = cdxi825m&cdxi643m;
wire cdxi3888m = cdxi825m&cdxi644m;
wire cdxi3889m = cdxi445m&cdxi913m;
wire cdxi3890m = cdxi582m&cdxi989m;
wire cdxi3891m = cdxi405m&cdxi1025m;
wire cdxi3892m = cdxi405m&cdxi1026m;
wire cdxi3893m = cdxi1013m&r33m;
wire cdxi3894m = cdxi977m&r34m;
wire cdxi3895m = cdxi1304m&r35m;
wire cdxi3896m = cdxi900m&r37m;
wire cdxi3897m = cdxi861m&r38m;
wire cdxi3898m = cdxi822m&r40m;
wire cdxi3899m = cdxi1014m&r43m;
wire cdxi3900m = cdxi978m&r44m;
wire cdxi3901m = cdxi1233m&r45m;
wire cdxi3902m = cdxi901m&r47m;
wire cdxi3903m = cdxi862m&r48m;
wire cdxi3904m = cdxi823m&r50m;
wire cdxi3905m = cdxi902m&r53m;
wire cdxi3906m = cdxi863m&r54m;
wire cdxi3907m = cdxi824m&r56m;
wire cdxi3908m = cdxi825m&r59m;
wire cdxi3909m = cdxi638m&r63m;
wire cdxi3910m = cdxi466m&r64m;
wire cdxi3911m = cdxi445m&r65m;
wire cdxi3912m = cdxi601m&r67m;
wire cdxi3913m = cdxi582m&r68m;
wire cdxi3914m = cdxi405m&r70m;
wire cdxi3915m = cdxi384m&r73m;
wire cdxi3916m = cdxi524m&r74m;
wire cdxi3917m = cdxi504m&r76m;
wire cdxi3918m = cdxi361m&r79m;
wire cdxi3919m = cdxi385m&r83m;
wire cdxi3920m = cdxi446m&r84m;
wire cdxi3921m = cdxi406m&r86m;
wire cdxi3922m = cdxi362m&r89m;
wire cdxi3923m = cdxi363m&r93m;
wire cdxi3924m = cdxi218m&r98m;
wire cdxi3925m = cdxi240m&r99m;
wire cdxi3926m = cdxi196m&r101m;
wire cdxi3927m = cdxi184m&r104m;
wire cdxi3928m = cdxi219m&r108m;
wire cdxi3929m = cdxi185m&r113m;
wire cdxi3930m = (cdxi3865m ^ cdxi3868m ^ cdxi3869m ^ cdxi3870m ^ cdxi3871m ^ cdxi3872m ^ cdxi3873m ^ cdxi3874m ^ cdxi3875m ^ cdxi3876m ^ cdxi3877m ^ cdxi3878m ^ cdxi3879m ^ cdxi3880m ^ cdxi3881m ^ cdxi3882m ^ cdxi3883m ^ cdxi3884m ^ cdxi3885m ^ cdxi3886m ^ cdxi3887m ^ cdxi3888m ^ cdxi3889m ^ cdxi3890m ^ cdxi3891m ^ cdxi3892m ^ cdxi3893m ^ cdxi3894m ^ cdxi3895m ^ cdxi3896m ^ cdxi3897m ^ cdxi3898m ^ cdxi3899m ^ cdxi3900m ^ cdxi3901m ^ cdxi3902m ^ cdxi3903m ^ cdxi3904m ^ cdxi3905m ^ cdxi3906m ^ cdxi3907m ^ cdxi3908m ^ cdxi3909m ^ cdxi3910m ^ cdxi3911m ^ cdxi3912m ^ cdxi3913m ^ cdxi3914m ^ cdxi3915m ^ cdxi3916m ^ cdxi3917m ^ cdxi3918m ^ cdxi3919m ^ cdxi3920m ^ cdxi3921m ^ cdxi3922m ^ cdxi3923m ^ cdxi3924m ^ cdxi3925m ^ cdxi3926m ^ cdxi3927m ^ cdxi3928m ^ cdxi3929m);
wire cdxi3931m = a0&cdxi3930m;
wire cdxi3932m = (reg_0_127);
wire cdxi3933m = reg_0_2&cdxi2290m;
wire cdxi3934m = reg_0_1&cdxi3833m;
wire cdxi3935m = reg_0_1&cdxi3834m;
wire cdxi3936m = reg_0_1&cdxi3835m;
wire cdxi3937m = reg_0_1&cdxi3836m;
wire cdxi3938m = reg_0_1&cdxi3837m;
wire cdxi3939m = reg_0_3&cdxi2086m;
wire cdxi3940m = reg_0_2&cdxi2295m;
wire cdxi3941m = reg_0_2&cdxi2296m;
wire cdxi3942m = reg_0_2&cdxi2297m;
wire cdxi3943m = reg_0_2&cdxi2298m;
wire cdxi3944m = reg_0_1&cdxi3838m;
wire cdxi3945m = reg_0_1&cdxi3839m;
wire cdxi3946m = reg_0_1&cdxi3840m;
wire cdxi3947m = reg_0_1&cdxi3841m;
wire cdxi3948m = reg_0_1&cdxi3842m;
wire cdxi3949m = reg_0_1&cdxi3843m;
wire cdxi3950m = reg_0_1&cdxi3844m;
wire cdxi3951m = reg_0_1&cdxi3845m;
wire cdxi3952m = reg_0_1&cdxi3846m;
wire cdxi3953m = reg_0_1&cdxi3847m;
wire cdxi3954m = reg_0_4&cdxi1956m;
wire cdxi3955m = reg_0_3&cdxi2096m;
wire cdxi3956m = reg_0_3&cdxi2097m;
wire cdxi3957m = reg_0_3&cdxi2098m;
wire cdxi3958m = reg_0_2&cdxi2305m;
wire cdxi3959m = reg_0_2&cdxi2306m;
wire cdxi3960m = reg_0_2&cdxi2307m;
wire cdxi3961m = reg_0_2&cdxi2308m;
wire cdxi3962m = reg_0_2&cdxi2309m;
wire cdxi3963m = reg_0_2&cdxi2310m;
wire cdxi3964m = reg_0_1&cdxi3848m;
wire cdxi3965m = reg_0_1&cdxi3849m;
wire cdxi3966m = reg_0_1&cdxi3850m;
wire cdxi3967m = reg_0_1&cdxi3851m;
wire cdxi3968m = reg_0_1&cdxi3852m;
wire cdxi3969m = reg_0_1&cdxi3853m;
wire cdxi3970m = reg_0_1&cdxi3854m;
wire cdxi3971m = reg_0_1&cdxi3855m;
wire cdxi3972m = reg_0_1&cdxi3856m;
wire cdxi3973m = reg_0_1&cdxi3857m;
wire cdxi3974m = reg_0_5&cdxi1896m;
wire cdxi3975m = reg_0_4&cdxi1966m;
wire cdxi3976m = reg_0_4&cdxi1967m;
wire cdxi3977m = reg_0_3&cdxi2106m;
wire cdxi3978m = reg_0_3&cdxi2107m;
wire cdxi3979m = reg_0_3&cdxi2108m;
wire cdxi3980m = reg_0_2&cdxi2315m;
wire cdxi3981m = reg_0_2&cdxi2316m;
wire cdxi3982m = reg_0_2&cdxi2317m;
wire cdxi3983m = reg_0_2&cdxi2318m;
wire cdxi3984m = reg_0_1&cdxi3858m;
wire cdxi3985m = reg_0_1&cdxi3859m;
wire cdxi3986m = reg_0_1&cdxi3860m;
wire cdxi3987m = reg_0_1&cdxi3861m;
wire cdxi3988m = reg_0_1&cdxi3862m;
wire cdxi3989m = reg_0_6&cdxi1800m;
wire cdxi3990m = reg_0_5&cdxi1870m;
wire cdxi3991m = reg_0_4&cdxi1940m;
wire cdxi3992m = reg_0_3&cdxi2080m;
wire cdxi3993m = reg_0_2&cdxi2289m;
wire cdxi3994m = reg_0_1&cdxi3832m;
wire cdxi3995m = (cdxi3933m ^ cdxi3934m ^ cdxi3935m ^ cdxi3936m ^ cdxi3937m ^ cdxi3938m ^ cdxi3939m ^ cdxi3940m ^ cdxi3941m ^ cdxi3942m ^ cdxi3943m ^ cdxi3944m ^ cdxi3945m ^ cdxi3946m ^ cdxi3947m ^ cdxi3948m ^ cdxi3949m ^ cdxi3950m ^ cdxi3951m ^ cdxi3952m ^ cdxi3953m ^ cdxi3954m ^ cdxi3955m ^ cdxi3956m ^ cdxi3957m ^ cdxi3958m ^ cdxi3959m ^ cdxi3960m ^ cdxi3961m ^ cdxi3962m ^ cdxi3963m ^ cdxi3964m ^ cdxi3965m ^ cdxi3966m ^ cdxi3967m ^ cdxi3968m ^ cdxi3969m ^ cdxi3970m ^ cdxi3971m ^ cdxi3972m ^ cdxi3973m ^ cdxi3974m ^ cdxi3975m ^ cdxi3976m ^ cdxi3977m ^ cdxi3978m ^ cdxi3979m ^ cdxi3980m ^ cdxi3981m ^ cdxi3982m ^ cdxi3983m ^ cdxi3984m ^ cdxi3985m ^ cdxi3986m ^ cdxi3987m ^ cdxi3988m ^ cdxi3989m ^ cdxi3990m ^ cdxi3991m ^ cdxi3992m ^ cdxi3993m ^ cdxi3994m ^ cdxi3932m);
wire cdxi3996m = reg_0_0&cdxi3995m;
wire cdxi3997m = cdxi1761m&cdxi657m ^ r125m;
wire cdxi3998m = cdxi361m&cdxi1232m;
wire cdxi3999m = cdxi2256m&cdxi271m;
wire cdxi4000m = cdxi2045m&cdxi230m;
wire cdxi4001m = cdxi361m&cdxi1727m;
wire cdxi4002m = cdxi361m&cdxi1728m;
wire cdxi4003m = cdxi361m&cdxi1729m;
wire cdxi4004m = cdxi361m&cdxi1730m;
wire cdxi4005m = cdxi445m&cdxi1449m;
wire cdxi4006m = cdxi1374m&cdxi567m;
wire cdxi4007m = cdxi2527m&r15m;
wire cdxi4008m = cdxi2323m&r16m;
wire cdxi4009m = cdxi2256m&r17m;
wire cdxi4010m = cdxi524m&cdxi1657m;
wire cdxi4011m = cdxi977m&cdxi623m;
wire cdxi4012m = cdxi2459m&r20m;
wire cdxi4013m = cdxi2045m&r21m;
wire cdxi4014m = cdxi361m&cdxi1731m;
wire cdxi4015m = cdxi361m&cdxi1732m;
wire cdxi4016m = cdxi361m&cdxi1733m;
wire cdxi4017m = cdxi361m&cdxi1734m;
wire cdxi4018m = cdxi361m&cdxi1735m;
wire cdxi4019m = cdxi361m&cdxi1736m;
wire cdxi4020m = cdxi638m&cdxi1350m;
wire cdxi4021m = cdxi1268m&r44m;
wire cdxi4022m = cdxi1232m&r45m;
wire cdxi4023m = cdxi445m&cdxi1456m;
wire cdxi4024m = cdxi1196m&r47m;
wire cdxi4025m = cdxi1160m&r48m;
wire cdxi4026m = cdxi1374m&r49m;
wire cdxi4027m = cdxi1123m&r50m;
wire cdxi4028m = cdxi1088m&r51m;
wire cdxi4029m = cdxi1303m&r52m;
wire cdxi4030m = cdxi1050m&r53m;
wire cdxi4031m = cdxi1410m&r54m;
wire cdxi4032m = cdxi1013m&r55m;
wire cdxi4033m = cdxi1339m&r56m;
wire cdxi4034m = cdxi977m&r57m;
wire cdxi4035m = cdxi1304m&r58m;
wire cdxi4036m = cdxi938m&r59m;
wire cdxi4037m = cdxi900m&r60m;
wire cdxi4038m = cdxi861m&r61m;
wire cdxi4039m = cdxi822m&r62m;
wire cdxi4040m = cdxi657m&r83m;
wire cdxi4041m = cdxi485m&r84m;
wire cdxi4042m = cdxi638m&r85m;
wire cdxi4043m = cdxi562m&r86m;
wire cdxi4044m = cdxi466m&r87m;
wire cdxi4045m = cdxi445m&r88m;
wire cdxi4046m = cdxi425m&r89m;
wire cdxi4047m = cdxi601m&r90m;
wire cdxi4048m = cdxi582m&r91m;
wire cdxi4049m = cdxi405m&r92m;
wire cdxi4050m = cdxi563m&r93m;
wire cdxi4051m = cdxi384m&r94m;
wire cdxi4052m = cdxi524m&r95m;
wire cdxi4053m = cdxi504m&r96m;
wire cdxi4054m = cdxi361m&r97m;
wire cdxi4055m = cdxi207m&r113m;
wire cdxi4056m = cdxi218m&r114m;
wire cdxi4057m = cdxi240m&r115m;
wire cdxi4058m = cdxi196m&r116m;
wire cdxi4059m = cdxi184m&r117m;
wire cdxi4060m = cdxi219m&r118m;
wire cdxi4061m = (cdxi3997m ^ cdxi3999m ^ cdxi4000m ^ cdxi4001m ^ cdxi4002m ^ cdxi4003m ^ cdxi4004m ^ cdxi4005m ^ cdxi4006m ^ cdxi4007m ^ cdxi4008m ^ cdxi4009m ^ cdxi4010m ^ cdxi4011m ^ cdxi4012m ^ cdxi4013m ^ cdxi4014m ^ cdxi4015m ^ cdxi4016m ^ cdxi4017m ^ cdxi4018m ^ cdxi4019m ^ cdxi4020m ^ cdxi4021m ^ cdxi4022m ^ cdxi4023m ^ cdxi4024m ^ cdxi4025m ^ cdxi4026m ^ cdxi4027m ^ cdxi4028m ^ cdxi4029m ^ cdxi4030m ^ cdxi4031m ^ cdxi4032m ^ cdxi4033m ^ cdxi4034m ^ cdxi4035m ^ cdxi4036m ^ cdxi4037m ^ cdxi4038m ^ cdxi4039m ^ cdxi4040m ^ cdxi4041m ^ cdxi4042m ^ cdxi4043m ^ cdxi4044m ^ cdxi4045m ^ cdxi4046m ^ cdxi4047m ^ cdxi4048m ^ cdxi4049m ^ cdxi4050m ^ cdxi4051m ^ cdxi4052m ^ cdxi4053m ^ cdxi4054m ^ cdxi4055m ^ cdxi4056m ^ cdxi4057m ^ cdxi4058m ^ cdxi4059m ^ cdxi4060m);
wire cdxi4062m = a0&cdxi4061m;
wire cdxi4063m = (reg_0_133);
wire cdxi4064m = reg_0_3&cdxi2628m;
wire cdxi4065m = reg_0_2&cdxi2695m;
wire cdxi4066m = reg_0_2&cdxi2696m;
wire cdxi4067m = reg_0_2&cdxi2697m;
wire cdxi4068m = reg_0_2&cdxi2698m;
wire cdxi4069m = reg_0_2&cdxi2699m;
wire cdxi4070m = reg_0_4&cdxi2770m;
wire cdxi4071m = reg_0_3&cdxi2633m;
wire cdxi4072m = reg_0_3&cdxi2634m;
wire cdxi4073m = reg_0_3&cdxi2635m;
wire cdxi4074m = reg_0_3&cdxi2636m;
wire cdxi4075m = reg_0_2&cdxi2700m;
wire cdxi4076m = reg_0_2&cdxi2701m;
wire cdxi4077m = reg_0_2&cdxi2702m;
wire cdxi4078m = reg_0_2&cdxi2703m;
wire cdxi4079m = reg_0_2&cdxi2704m;
wire cdxi4080m = reg_0_2&cdxi2705m;
wire cdxi4081m = reg_0_2&cdxi2706m;
wire cdxi4082m = reg_0_2&cdxi2707m;
wire cdxi4083m = reg_0_2&cdxi2708m;
wire cdxi4084m = reg_0_2&cdxi2709m;
wire cdxi4085m = reg_0_5&cdxi2577m;
wire cdxi4086m = reg_0_4&cdxi2780m;
wire cdxi4087m = reg_0_4&cdxi2781m;
wire cdxi4088m = reg_0_4&cdxi2782m;
wire cdxi4089m = reg_0_3&cdxi2643m;
wire cdxi4090m = reg_0_3&cdxi2644m;
wire cdxi4091m = reg_0_3&cdxi2645m;
wire cdxi4092m = reg_0_3&cdxi2646m;
wire cdxi4093m = reg_0_3&cdxi2647m;
wire cdxi4094m = reg_0_3&cdxi2648m;
wire cdxi4095m = reg_0_2&cdxi2710m;
wire cdxi4096m = reg_0_2&cdxi2711m;
wire cdxi4097m = reg_0_2&cdxi2712m;
wire cdxi4098m = reg_0_2&cdxi2713m;
wire cdxi4099m = reg_0_2&cdxi2714m;
wire cdxi4100m = reg_0_2&cdxi2715m;
wire cdxi4101m = reg_0_2&cdxi2716m;
wire cdxi4102m = reg_0_2&cdxi2717m;
wire cdxi4103m = reg_0_2&cdxi2718m;
wire cdxi4104m = reg_0_2&cdxi2719m;
wire cdxi4105m = reg_0_6&cdxi2519m;
wire cdxi4106m = reg_0_5&cdxi2587m;
wire cdxi4107m = reg_0_5&cdxi2588m;
wire cdxi4108m = reg_0_4&cdxi2790m;
wire cdxi4109m = reg_0_4&cdxi2791m;
wire cdxi4110m = reg_0_4&cdxi2792m;
wire cdxi4111m = reg_0_3&cdxi2653m;
wire cdxi4112m = reg_0_3&cdxi2654m;
wire cdxi4113m = reg_0_3&cdxi2655m;
wire cdxi4114m = reg_0_3&cdxi2656m;
wire cdxi4115m = reg_0_2&cdxi2720m;
wire cdxi4116m = reg_0_2&cdxi2721m;
wire cdxi4117m = reg_0_2&cdxi2722m;
wire cdxi4118m = reg_0_2&cdxi2723m;
wire cdxi4119m = reg_0_2&cdxi2724m;
wire cdxi4120m = reg_0_7&cdxi3832m;
wire cdxi4121m = reg_0_6&cdxi2493m;
wire cdxi4122m = reg_0_5&cdxi2561m;
wire cdxi4123m = reg_0_4&cdxi2764m;
wire cdxi4124m = reg_0_3&cdxi2627m;
wire cdxi4125m = reg_0_2&cdxi2694m;
wire cdxi4126m = (cdxi4064m ^ cdxi4065m ^ cdxi4066m ^ cdxi4067m ^ cdxi4068m ^ cdxi4069m ^ cdxi4070m ^ cdxi4071m ^ cdxi4072m ^ cdxi4073m ^ cdxi4074m ^ cdxi4075m ^ cdxi4076m ^ cdxi4077m ^ cdxi4078m ^ cdxi4079m ^ cdxi4080m ^ cdxi4081m ^ cdxi4082m ^ cdxi4083m ^ cdxi4084m ^ cdxi4085m ^ cdxi4086m ^ cdxi4087m ^ cdxi4088m ^ cdxi4089m ^ cdxi4090m ^ cdxi4091m ^ cdxi4092m ^ cdxi4093m ^ cdxi4094m ^ cdxi4095m ^ cdxi4096m ^ cdxi4097m ^ cdxi4098m ^ cdxi4099m ^ cdxi4100m ^ cdxi4101m ^ cdxi4102m ^ cdxi4103m ^ cdxi4104m ^ cdxi4105m ^ cdxi4106m ^ cdxi4107m ^ cdxi4108m ^ cdxi4109m ^ cdxi4110m ^ cdxi4111m ^ cdxi4112m ^ cdxi4113m ^ cdxi4114m ^ cdxi4115m ^ cdxi4116m ^ cdxi4117m ^ cdxi4118m ^ cdxi4119m ^ cdxi4120m ^ cdxi4121m ^ cdxi4122m ^ cdxi4123m ^ cdxi4124m ^ cdxi4125m ^ cdxi4063m);
wire cdxi4127m = reg_0_0&cdxi4126m;
wire cdxi4128m = cdxi185m ^ cdxi184m ^ cdxi240m ^ cdxi218m;
wire cdxi4129m = cdxi185m&cdxi152m;
wire cdxi4130m = reg_0_1&cdxi155m;
wire cdxi4131m = cdxi219m&cdxi168m;
wire cdxi4132m = reg_0_2&cdxi171m;
wire cdxi4133m = cdxi184m&cdxi168m;
wire cdxi4134m = reg_0_3&cdxi171m;
wire cdxi4135m = cdxi361m ^ r13m;
wire cdxi4136m = cdxi184m&r1m;
wire cdxi4137m = cdxi219m&r2m;
wire cdxi4138m = (cdxi4135m ^ cdxi4136m ^ cdxi4137m);
wire cdxi4139m = cdxi185m&cdxi4138m;
wire cdxi4140m = reg_0_3&cdxi136m;
wire cdxi4141m = reg_0_2&cdxi142m;
wire cdxi4142m = (cdxi4140m ^ cdxi4141m ^ cdxi373m);
wire cdxi4143m = reg_0_1&cdxi4142m;
wire cdxi4144m = cdxi185m&cdxi222m;
wire cdxi4145m = reg_0_1&cdxi227m;
wire cdxi4146m = cdxi185m&cdxi313m;
wire cdxi4147m = reg_0_1&cdxi318m;
wire cdxi4148m = cdxi185m&cdxi263m;
wire cdxi4149m = reg_0_1&cdxi268m;
wire cdxi4150m = cdxi185m&cdxi339m;
wire cdxi4151m = reg_0_1&cdxi344m;
wire cdxi4152m = cdxi196m&cdxi339m;
wire cdxi4153m = reg_0_4&cdxi344m;
wire cdxi4154m = cdxi1014m ^ r40m;
wire cdxi4155m = cdxi638m&r0m;
wire cdxi4156m = cdxi185m&cdxi251m;
wire cdxi4157m = cdxi185m&cdxi252m;
wire cdxi4158m = cdxi218m&r10m;
wire cdxi4159m = cdxi240m&r11m;
wire cdxi4160m = cdxi185m&r25m;
wire cdxi4161m = (cdxi4154m ^ cdxi4155m ^ cdxi4156m ^ cdxi4157m ^ cdxi4158m ^ cdxi4159m ^ cdxi4160m);
wire cdxi4162m = a0&cdxi4161m;
wire cdxi4163m = reg_0_5&reg_0_6&cdxi130m;
wire cdxi4164m = reg_0_1&cdxi256m;
wire cdxi4165m = reg_0_1&cdxi257m;
wire cdxi4166m = reg_0_6&cdxi455m;
wire cdxi4167m = reg_0_5&cdxi394m;
wire cdxi4168m = reg_0_1&cdxi255m;
wire cdxi4169m = (cdxi4163m ^ cdxi4164m ^ cdxi4165m ^ cdxi4166m ^ cdxi4167m ^ cdxi4168m ^ cdxi1031m);
wire cdxi4170m = reg_0_0&cdxi4169m;
wire cdxi4171m = cdxi1051m ^ r42m;
wire cdxi4172m = cdxi218m&cdxi208m;
wire cdxi4173m = cdxi185m&cdxi337m;
wire cdxi4174m = cdxi185m&cdxi338m;
wire cdxi4175m = cdxi207m&r11m;
wire cdxi4176m = cdxi218m&r12m;
wire cdxi4177m = cdxi185m&r27m;
wire cdxi4178m = (cdxi4171m ^ cdxi4172m ^ cdxi4173m ^ cdxi4174m ^ cdxi4175m ^ cdxi4176m ^ cdxi4177m);
wire cdxi4179m = a0&cdxi4178m;
wire cdxi4180m = reg_0_6&cdxi213m;
wire cdxi4181m = reg_0_1&cdxi342m;
wire cdxi4182m = reg_0_1&cdxi343m;
wire cdxi4183m = reg_0_7&cdxi394m;
wire cdxi4184m = reg_0_6&cdxi212m;
wire cdxi4185m = reg_0_1&cdxi341m;
wire cdxi4186m = (cdxi4180m ^ cdxi4181m ^ cdxi4182m ^ cdxi4183m ^ cdxi4184m ^ cdxi4185m ^ cdxi1068m);
wire cdxi4187m = reg_0_0&cdxi4186m;
wire cdxi4188m = a0&cdxi682m;
wire cdxi4189m = reg_0_0&cdxi691m;
wire cdxi4190m = a0&cdxi722m;
wire cdxi4191m = reg_0_0&cdxi731m;
wire cdxi4192m = cdxi185m&cdxi3568m;
wire cdxi4193m = reg_0_1&cdxi3576m;
wire cdxi4194m = cdxi185m&cdxi808m;
wire cdxi4195m = reg_0_1&cdxi817m;
wire cdxi4196m = cdxi2046m ^ r79m;
wire cdxi4197m = cdxi1479m&r0m;
wire cdxi4198m = cdxi446m&cdxi301m;
wire cdxi4199m = cdxi406m&cdxi251m;
wire cdxi4200m = cdxi406m&cdxi252m;
wire cdxi4201m = cdxi240m&cdxi470m;
wire cdxi4202m = cdxi466m&r10m;
wire cdxi4203m = cdxi445m&r11m;
wire cdxi4204m = cdxi385m&r22m;
wire cdxi4205m = cdxi446m&r23m;
wire cdxi4206m = cdxi406m&r25m;
wire cdxi4207m = cdxi218m&r37m;
wire cdxi4208m = cdxi240m&r38m;
wire cdxi4209m = cdxi196m&r40m;
wire cdxi4210m = cdxi185m&r59m;
wire cdxi4211m = (cdxi4196m ^ cdxi4197m ^ cdxi4198m ^ cdxi4199m ^ cdxi4200m ^ cdxi4201m ^ cdxi4202m ^ cdxi4203m ^ cdxi4204m ^ cdxi4205m ^ cdxi4206m ^ cdxi4207m ^ cdxi4208m ^ cdxi4209m ^ cdxi4210m);
wire cdxi4212m = a0&cdxi4211m;
wire cdxi4213m = reg_0_4&cdxi4163m;
wire cdxi4214m = reg_0_1&cdxi648m;
wire cdxi4215m = reg_0_1&cdxi649m;
wire cdxi4216m = reg_0_1&cdxi650m;
wire cdxi4217m = reg_0_5&cdxi479m;
wire cdxi4218m = reg_0_4&cdxi4166m;
wire cdxi4219m = reg_0_4&cdxi4167m;
wire cdxi4220m = reg_0_1&cdxi651m;
wire cdxi4221m = reg_0_1&cdxi652m;
wire cdxi4222m = reg_0_1&cdxi653m;
wire cdxi4223m = reg_0_6&cdxi456m;
wire cdxi4224m = reg_0_5&cdxi475m;
wire cdxi4225m = reg_0_4&cdxi1031m;
wire cdxi4226m = reg_0_1&cdxi647m;
wire cdxi4227m = (cdxi4213m ^ cdxi4214m ^ cdxi4215m ^ cdxi4216m ^ cdxi4217m ^ cdxi4218m ^ cdxi4219m ^ cdxi4220m ^ cdxi4221m ^ cdxi4222m ^ cdxi4223m ^ cdxi4224m ^ cdxi4225m ^ cdxi4226m ^ cdxi2079m);
wire cdxi4228m = reg_0_0&cdxi4227m;
wire cdxi4229m = a0&cdxi1633m;
wire cdxi4230m = reg_0_0&cdxi1650m;
wire cdxi4231m = cdxi185m&cdxi1494m;
wire cdxi4232m = reg_0_1&cdxi1511m;
wire cdxi4233m = cdxi185m&cdxi3665m;
wire cdxi4234m = reg_0_1&cdxi3681m;
wire cdxi4235m = cdxi185m&cdxi1701m;
wire cdxi4236m = reg_0_1&cdxi1718m;
wire cdxi4237m = cdxi2941m ^ r111m;
wire cdxi4238m = cdxi1374m&cdxi208m;
wire cdxi4239m = cdxi1014m&cdxi230m;
wire cdxi4240m = cdxi362m&cdxi658m;
wire cdxi4241m = cdxi362m&cdxi659m;
wire cdxi4242m = cdxi362m&cdxi660m;
wire cdxi4243m = cdxi638m&cdxi430m;
wire cdxi4244m = cdxi601m&cdxi489m;
wire cdxi4245m = cdxi1160m&r11m;
wire cdxi4246m = cdxi1374m&r12m;
wire cdxi4247m = cdxi385m&cdxi623m;
wire cdxi4248m = cdxi1161m&r20m;
wire cdxi4249m = cdxi1014m&r21m;
wire cdxi4250m = cdxi362m&cdxi661m;
wire cdxi4251m = cdxi362m&cdxi662m;
wire cdxi4252m = cdxi362m&cdxi663m;
wire cdxi4253m = cdxi657m&r34m;
wire cdxi4254m = cdxi485m&r35m;
wire cdxi4255m = cdxi638m&r36m;
wire cdxi4256m = cdxi425m&r40m;
wire cdxi4257m = cdxi601m&r41m;
wire cdxi4258m = cdxi582m&r42m;
wire cdxi4259m = cdxi426m&r56m;
wire cdxi4260m = cdxi385m&r57m;
wire cdxi4261m = cdxi446m&r58m;
wire cdxi4262m = cdxi362m&r62m;
wire cdxi4263m = cdxi207m&r76m;
wire cdxi4264m = cdxi218m&r77m;
wire cdxi4265m = cdxi240m&r78m;
wire cdxi4266m = cdxi184m&r82m;
wire cdxi4267m = cdxi185m&r96m;
wire cdxi4268m = (cdxi4237m ^ cdxi4238m ^ cdxi4239m ^ cdxi4240m ^ cdxi4241m ^ cdxi4242m ^ cdxi4243m ^ cdxi4244m ^ cdxi4245m ^ cdxi4246m ^ cdxi4247m ^ cdxi4248m ^ cdxi4249m ^ cdxi4250m ^ cdxi4251m ^ cdxi4252m ^ cdxi4253m ^ cdxi4254m ^ cdxi4255m ^ cdxi4256m ^ cdxi4257m ^ cdxi4258m ^ cdxi4259m ^ cdxi4260m ^ cdxi4261m ^ cdxi4262m ^ cdxi4263m ^ cdxi4264m ^ cdxi4265m ^ cdxi4266m ^ cdxi4267m);
wire cdxi4269m = a0&cdxi4268m;
wire cdxi4270m = reg_0_3&cdxi3634m;
wire cdxi4271m = reg_0_1&cdxi1566m;
wire cdxi4272m = reg_0_1&cdxi1567m;
wire cdxi4273m = reg_0_1&cdxi1568m;
wire cdxi4274m = reg_0_1&cdxi1569m;
wire cdxi4275m = reg_0_5&cdxi1219m;
wire cdxi4276m = reg_0_3&cdxi3638m;
wire cdxi4277m = reg_0_3&cdxi3639m;
wire cdxi4278m = reg_0_3&cdxi3640m;
wire cdxi4279m = reg_0_1&cdxi1570m;
wire cdxi4280m = reg_0_1&cdxi1571m;
wire cdxi4281m = reg_0_1&cdxi1572m;
wire cdxi4282m = reg_0_1&cdxi1573m;
wire cdxi4283m = reg_0_1&cdxi1574m;
wire cdxi4284m = reg_0_1&cdxi1575m;
wire cdxi4285m = reg_0_6&cdxi1189m;
wire cdxi4286m = reg_0_5&cdxi1225m;
wire cdxi4287m = reg_0_5&cdxi1226m;
wire cdxi4288m = reg_0_3&cdxi3644m;
wire cdxi4289m = reg_0_3&cdxi3645m;
wire cdxi4290m = reg_0_3&cdxi3646m;
wire cdxi4291m = reg_0_1&cdxi1576m;
wire cdxi4292m = reg_0_1&cdxi1577m;
wire cdxi4293m = reg_0_1&cdxi1578m;
wire cdxi4294m = reg_0_1&cdxi1579m;
wire cdxi4295m = reg_0_7&cdxi1939m;
wire cdxi4296m = reg_0_6&cdxi1178m;
wire cdxi4297m = reg_0_5&cdxi1214m;
wire cdxi4298m = reg_0_3&cdxi2220m;
wire cdxi4299m = reg_0_1&cdxi1565m;
wire cdxi4300m = (cdxi4270m ^ cdxi4271m ^ cdxi4272m ^ cdxi4273m ^ cdxi4274m ^ cdxi4275m ^ cdxi4276m ^ cdxi4277m ^ cdxi4278m ^ cdxi4279m ^ cdxi4280m ^ cdxi4281m ^ cdxi4282m ^ cdxi4283m ^ cdxi4284m ^ cdxi4285m ^ cdxi4286m ^ cdxi4287m ^ cdxi4288m ^ cdxi4289m ^ cdxi4290m ^ cdxi4291m ^ cdxi4292m ^ cdxi4293m ^ cdxi4294m ^ cdxi4295m ^ cdxi4296m ^ cdxi4297m ^ cdxi4298m ^ cdxi4299m ^ cdxi3009m);
wire cdxi4301m = reg_0_0&cdxi4300m;
wire cdxi4302m = cdxi185m&cdxi2625m;
wire cdxi4303m = reg_0_1&cdxi2658m;
wire cdxi4304m = cdxi219m&cdxi2692m;
wire cdxi4305m = reg_0_2&cdxi2725m;
wire cdxi4306m = cdxi825m&cdxi1232m ^ r120m;
wire cdxi4307m = cdxi361m&cdxi1234m;
wire cdxi4308m = cdxi362m&cdxi1514m;
wire cdxi4309m = cdxi363m&cdxi1619m;
wire cdxi4310m = cdxi825m&cdxi802m;
wire cdxi4311m = cdxi825m&cdxi803m;
wire cdxi4312m = cdxi825m&cdxi804m;
wire cdxi4313m = cdxi2323m&r7m;
wire cdxi4314m = cdxi1304m&cdxi430m;
wire cdxi4315m = cdxi361m&cdxi1238m;
wire cdxi4316m = cdxi822m&cdxi489m;
wire cdxi4317m = cdxi361m&cdxi1240m;
wire cdxi4318m = cdxi406m&cdxi1415m;
wire cdxi4319m = cdxi362m&cdxi1518m;
wire cdxi4320m = cdxi362m&cdxi1519m;
wire cdxi4321m = cdxi362m&cdxi1520m;
wire cdxi4322m = cdxi363m&cdxi1623m;
wire cdxi4323m = cdxi363m&cdxi1624m;
wire cdxi4324m = cdxi363m&cdxi1625m;
wire cdxi4325m = cdxi825m&cdxi805m;
wire cdxi4326m = cdxi825m&cdxi806m;
wire cdxi4327m = cdxi825m&cdxi807m;
wire cdxi4328m = cdxi445m&cdxi951m;
wire cdxi4329m = cdxi1160m&r29m;
wire cdxi4330m = cdxi1123m&r30m;
wire cdxi4331m = cdxi1303m&r32m;
wire cdxi4332m = cdxi1410m&r33m;
wire cdxi4333m = cdxi504m&cdxi1172m;
wire cdxi4334m = cdxi1304m&r36m;
wire cdxi4335m = cdxi938m&r37m;
wire cdxi4336m = cdxi861m&r39m;
wire cdxi4337m = cdxi822m&r41m;
wire cdxi4338m = cdxi1161m&r43m;
wire cdxi4339m = cdxi1124m&r44m;
wire cdxi4340m = cdxi1233m&r46m;
wire cdxi4341m = cdxi939m&r47m;
wire cdxi4342m = cdxi862m&r49m;
wire cdxi4343m = cdxi823m&r51m;
wire cdxi4344m = cdxi940m&r53m;
wire cdxi4345m = cdxi863m&r55m;
wire cdxi4346m = cdxi824m&r57m;
wire cdxi4347m = cdxi825m&r60m;
wire cdxi4348m = cdxi485m&r63m;
wire cdxi4349m = cdxi562m&r64m;
wire cdxi4350m = cdxi445m&r66m;
wire cdxi4351m = cdxi425m&r67m;
wire cdxi4352m = cdxi582m&r69m;
wire cdxi4353m = cdxi405m&r71m;
wire cdxi4354m = cdxi563m&r73m;
wire cdxi4355m = cdxi524m&r75m;
wire cdxi4356m = cdxi504m&r77m;
wire cdxi4357m = cdxi361m&r80m;
wire cdxi4358m = cdxi426m&r83m;
wire cdxi4359m = cdxi446m&r85m;
wire cdxi4360m = cdxi406m&r87m;
wire cdxi4361m = cdxi362m&r90m;
wire cdxi4362m = cdxi363m&r94m;
wire cdxi4363m = cdxi207m&r98m;
wire cdxi4364m = cdxi240m&r100m;
wire cdxi4365m = cdxi196m&r102m;
wire cdxi4366m = cdxi184m&r105m;
wire cdxi4367m = cdxi219m&r109m;
wire cdxi4368m = cdxi185m&r114m;
wire cdxi4369m = (cdxi4306m ^ cdxi4307m ^ cdxi4308m ^ cdxi4309m ^ cdxi4310m ^ cdxi4311m ^ cdxi4312m ^ cdxi4313m ^ cdxi4314m ^ cdxi4315m ^ cdxi4316m ^ cdxi4317m ^ cdxi4318m ^ cdxi4319m ^ cdxi4320m ^ cdxi4321m ^ cdxi4322m ^ cdxi4323m ^ cdxi4324m ^ cdxi4325m ^ cdxi4326m ^ cdxi4327m ^ cdxi4328m ^ cdxi4329m ^ cdxi4330m ^ cdxi4331m ^ cdxi4332m ^ cdxi4333m ^ cdxi4334m ^ cdxi4335m ^ cdxi4336m ^ cdxi4337m ^ cdxi4338m ^ cdxi4339m ^ cdxi4340m ^ cdxi4341m ^ cdxi4342m ^ cdxi4343m ^ cdxi4344m ^ cdxi4345m ^ cdxi4346m ^ cdxi4347m ^ cdxi4348m ^ cdxi4349m ^ cdxi4350m ^ cdxi4351m ^ cdxi4352m ^ cdxi4353m ^ cdxi4354m ^ cdxi4355m ^ cdxi4356m ^ cdxi4357m ^ cdxi4358m ^ cdxi4359m ^ cdxi4360m ^ cdxi4361m ^ cdxi4362m ^ cdxi4363m ^ cdxi4364m ^ cdxi4365m ^ cdxi4366m ^ cdxi4367m ^ cdxi4368m);
wire cdxi4370m = a0&cdxi4369m;
wire cdxi4371m = (reg_0_128);
wire cdxi4372m = reg_0_2&cdxi2359m;
wire cdxi4373m = reg_0_1&cdxi2494m;
wire cdxi4374m = reg_0_1&cdxi2495m;
wire cdxi4375m = reg_0_1&cdxi2496m;
wire cdxi4376m = reg_0_1&cdxi2497m;
wire cdxi4377m = reg_0_1&cdxi2498m;
wire cdxi4378m = reg_0_3&reg_0_4&reg_0_5&cdxi3451m;
wire cdxi4379m = reg_0_2&cdxi2364m;
wire cdxi4380m = reg_0_2&cdxi2365m;
wire cdxi4381m = reg_0_2&cdxi2366m;
wire cdxi4382m = reg_0_2&cdxi2367m;
wire cdxi4383m = reg_0_1&cdxi2499m;
wire cdxi4384m = reg_0_1&cdxi2500m;
wire cdxi4385m = reg_0_1&cdxi2501m;
wire cdxi4386m = reg_0_1&cdxi2502m;
wire cdxi4387m = reg_0_1&cdxi2503m;
wire cdxi4388m = reg_0_1&cdxi2504m;
wire cdxi4389m = reg_0_1&cdxi2505m;
wire cdxi4390m = reg_0_1&cdxi2506m;
wire cdxi4391m = reg_0_1&cdxi2507m;
wire cdxi4392m = reg_0_1&cdxi2508m;
wire cdxi4393m = reg_0_4&cdxi2027m;
wire cdxi4394m = reg_0_3&reg_0_5&cdxi3611m;
wire cdxi4395m = reg_0_3&reg_0_4&reg_0_7&cdxi880m;
wire cdxi4396m = reg_0_3&reg_0_4&reg_0_5&cdxi957m;
wire cdxi4397m = reg_0_2&cdxi2374m;
wire cdxi4398m = reg_0_2&cdxi2375m;
wire cdxi4399m = reg_0_2&cdxi2376m;
wire cdxi4400m = reg_0_2&cdxi2377m;
wire cdxi4401m = reg_0_2&cdxi2378m;
wire cdxi4402m = reg_0_2&cdxi2379m;
wire cdxi4403m = reg_0_1&cdxi2509m;
wire cdxi4404m = reg_0_1&cdxi2510m;
wire cdxi4405m = reg_0_1&cdxi2511m;
wire cdxi4406m = reg_0_1&cdxi2512m;
wire cdxi4407m = reg_0_1&cdxi2513m;
wire cdxi4408m = reg_0_1&cdxi2514m;
wire cdxi4409m = reg_0_1&cdxi2515m;
wire cdxi4410m = reg_0_1&cdxi2516m;
wire cdxi4411m = reg_0_1&cdxi2517m;
wire cdxi4412m = reg_0_1&cdxi2518m;
wire cdxi4413m = reg_0_5&reg_0_7&cdxi843m;
wire cdxi4414m = reg_0_4&cdxi2037m;
wire cdxi4415m = reg_0_4&cdxi2038m;
wire cdxi4416m = reg_0_3&reg_0_7&cdxi1798m;
wire cdxi4417m = reg_0_3&reg_0_5&cdxi2150m;
wire cdxi4418m = reg_0_3&reg_0_4&cdxi2010m;
wire cdxi4419m = reg_0_2&cdxi2384m;
wire cdxi4420m = reg_0_2&cdxi2385m;
wire cdxi4421m = reg_0_2&cdxi2386m;
wire cdxi4422m = reg_0_2&cdxi2387m;
wire cdxi4423m = reg_0_1&cdxi2519m;
wire cdxi4424m = reg_0_1&cdxi2520m;
wire cdxi4425m = reg_0_1&cdxi2521m;
wire cdxi4426m = reg_0_1&cdxi2522m;
wire cdxi4427m = reg_0_1&cdxi2523m;
wire cdxi4428m = reg_0_7&cdxi1800m;
wire cdxi4429m = reg_0_5&cdxi2871m;
wire cdxi4430m = reg_0_4&cdxi2011m;
wire cdxi4431m = reg_0_3&cdxi3144m;
wire cdxi4432m = reg_0_2&cdxi2358m;
wire cdxi4433m = reg_0_1&cdxi2493m;
wire cdxi4434m = (cdxi4372m ^ cdxi4373m ^ cdxi4374m ^ cdxi4375m ^ cdxi4376m ^ cdxi4377m ^ cdxi4378m ^ cdxi4379m ^ cdxi4380m ^ cdxi4381m ^ cdxi4382m ^ cdxi4383m ^ cdxi4384m ^ cdxi4385m ^ cdxi4386m ^ cdxi4387m ^ cdxi4388m ^ cdxi4389m ^ cdxi4390m ^ cdxi4391m ^ cdxi4392m ^ cdxi4393m ^ cdxi4394m ^ cdxi4395m ^ cdxi4396m ^ cdxi4397m ^ cdxi4398m ^ cdxi4399m ^ cdxi4400m ^ cdxi4401m ^ cdxi4402m ^ cdxi4403m ^ cdxi4404m ^ cdxi4405m ^ cdxi4406m ^ cdxi4407m ^ cdxi4408m ^ cdxi4409m ^ cdxi4410m ^ cdxi4411m ^ cdxi4412m ^ cdxi4413m ^ cdxi4414m ^ cdxi4415m ^ cdxi4416m ^ cdxi4417m ^ cdxi4418m ^ cdxi4419m ^ cdxi4420m ^ cdxi4421m ^ cdxi4422m ^ cdxi4423m ^ cdxi4424m ^ cdxi4425m ^ cdxi4426m ^ cdxi4427m ^ cdxi4428m ^ cdxi4429m ^ cdxi4430m ^ cdxi4431m ^ cdxi4432m ^ cdxi4433m ^ cdxi4371m);
wire cdxi4435m = reg_0_0&cdxi4434m;
wire cdxi4436m = cdxi185m&cdxi4061m;
wire cdxi4437m = reg_0_1&cdxi4126m;
wire cdxi4438m = 1&1 ^ cdxi185m ^ cdxi196m ^ cdxi218m ^ cdxi207m;
wire cdxi4439m = cdxi185m&cdxi232m;
wire cdxi4440m = reg_0_1&cdxi237m;
wire cdxi4441m = cdxi185m&cdxi243m;
wire cdxi4442m = reg_0_1&cdxi248m;
wire cdxi4443m = cdxi184m&cdxi339m;
wire cdxi4444m = reg_0_3&cdxi344m;
wire cdxi4445m = cdxi863m ^ r30m;
wire cdxi4446m = cdxi524m&r0m;
wire cdxi4447m = cdxi446m&r1m;
wire cdxi4448m = cdxi363m&r4m;
wire cdxi4449m = cdxi240m&r7m;
wire cdxi4450m = cdxi219m&r10m;
wire cdxi4451m = cdxi185m&r15m;
wire cdxi4452m = (cdxi4445m ^ cdxi4446m ^ cdxi4447m ^ cdxi4448m ^ cdxi4449m ^ cdxi4450m ^ cdxi4451m);
wire cdxi4453m = a0&cdxi4452m;
wire cdxi4454m = reg_0_2&cdxi3372m;
wire cdxi4455m = reg_0_1&cdxi3390m;
wire cdxi4456m = reg_0_1&cdxi3391m;
wire cdxi4457m = reg_0_5&cdxi372m;
wire cdxi4458m = reg_0_2&cdxi455m;
wire cdxi4459m = reg_0_1&cdxi533m;
wire cdxi4460m = (cdxi4454m ^ cdxi4455m ^ cdxi4456m ^ cdxi4457m ^ cdxi4458m ^ cdxi4459m ^ cdxi880m);
wire cdxi4461m = reg_0_0&cdxi4460m;
wire cdxi4462m = cdxi1976m ^ r71m;
wire cdxi4463m = cdxi219m&cdxi486m;
wire cdxi4464m = cdxi446m&cdxi271m;
wire cdxi4465m = cdxi363m&cdxi261m;
wire cdxi4466m = cdxi363m&cdxi262m;
wire cdxi4467m = cdxi485m&r7m;
wire cdxi4468m = cdxi219m&cdxi489m;
wire cdxi4469m = cdxi219m&cdxi490m;
wire cdxi4470m = cdxi426m&r15m;
wire cdxi4471m = cdxi446m&r17m;
wire cdxi4472m = cdxi363m&r26m;
wire cdxi4473m = cdxi207m&r30m;
wire cdxi4474m = cdxi240m&r32m;
wire cdxi4475m = cdxi219m&r41m;
wire cdxi4476m = cdxi185m&r51m;
wire cdxi4477m = (cdxi4462m ^ cdxi4463m ^ cdxi4464m ^ cdxi4465m ^ cdxi4466m ^ cdxi4467m ^ cdxi4468m ^ cdxi4469m ^ cdxi4470m ^ cdxi4471m ^ cdxi4472m ^ cdxi4473m ^ cdxi4474m ^ cdxi4475m ^ cdxi4476m);
wire cdxi4478m = a0&cdxi4477m;
wire cdxi4479m = reg_0_2&cdxi495m;
wire cdxi4480m = reg_0_1&cdxi743m;
wire cdxi4481m = reg_0_1&cdxi744m;
wire cdxi4482m = reg_0_1&cdxi745m;
wire cdxi4483m = reg_0_5&cdxi3451m;
wire cdxi4484m = reg_0_2&cdxi498m;
wire cdxi4485m = reg_0_2&cdxi499m;
wire cdxi4486m = reg_0_1&cdxi746m;
wire cdxi4487m = reg_0_1&cdxi747m;
wire cdxi4488m = reg_0_1&cdxi748m;
wire cdxi4489m = reg_0_7&cdxi880m;
wire cdxi4490m = reg_0_5&cdxi957m;
wire cdxi4491m = reg_0_2&cdxi494m;
wire cdxi4492m = reg_0_1&cdxi742m;
wire cdxi4493m = (cdxi4479m ^ cdxi4480m ^ cdxi4481m ^ cdxi4482m ^ cdxi4483m ^ cdxi4484m ^ cdxi4485m ^ cdxi4486m ^ cdxi4487m ^ cdxi4488m ^ cdxi4489m ^ cdxi4490m ^ cdxi4491m ^ cdxi4492m ^ cdxi2010m);
wire cdxi4494m = reg_0_0&cdxi4493m;
wire cdxi4495m = cdxi1762m ^ r73m;
wire cdxi4496m = cdxi1303m&r0m;
wire cdxi4497m = cdxi406m&cdxi311m;
wire cdxi4498m = cdxi362m&cdxi241m;
wire cdxi4499m = cdxi362m&cdxi242m;
wire cdxi4500m = cdxi445m&r8m;
wire cdxi4501m = cdxi184m&cdxi450m;
wire cdxi4502m = cdxi405m&r10m;
wire cdxi4503m = cdxi446m&r18m;
wire cdxi4504m = cdxi406m&r19m;
wire cdxi4505m = cdxi362m&r22m;
wire cdxi4506m = cdxi240m&r33m;
wire cdxi4507m = cdxi196m&r34m;
wire cdxi4508m = cdxi184m&r37m;
wire cdxi4509m = cdxi185m&r53m;
wire cdxi4510m = (cdxi4495m ^ cdxi4496m ^ cdxi4497m ^ cdxi4498m ^ cdxi4499m ^ cdxi4500m ^ cdxi4501m ^ cdxi4502m ^ cdxi4503m ^ cdxi4504m ^ cdxi4505m ^ cdxi4506m ^ cdxi4507m ^ cdxi4508m ^ cdxi4509m);
wire cdxi4511m = a0&cdxi4510m;
wire cdxi4512m = reg_0_3&cdxi457m;
wire cdxi4513m = reg_0_1&cdxi592m;
wire cdxi4514m = reg_0_1&cdxi593m;
wire cdxi4515m = reg_0_1&cdxi594m;
wire cdxi4516m = reg_0_4&cdxi3468m;
wire cdxi4517m = reg_0_3&cdxi460m;
wire cdxi4518m = reg_0_3&cdxi461m;
wire cdxi4519m = reg_0_1&cdxi595m;
wire cdxi4520m = reg_0_1&cdxi596m;
wire cdxi4521m = reg_0_1&cdxi597m;
wire cdxi4522m = reg_0_5&cdxi415m;
wire cdxi4523m = reg_0_4&cdxi881m;
wire cdxi4524m = reg_0_3&cdxi456m;
wire cdxi4525m = reg_0_1&cdxi591m;
wire cdxi4526m = (cdxi4512m ^ cdxi4513m ^ cdxi4514m ^ cdxi4515m ^ cdxi4516m ^ cdxi4517m ^ cdxi4518m ^ cdxi4519m ^ cdxi4520m ^ cdxi4521m ^ cdxi4522m ^ cdxi4523m ^ cdxi4524m ^ cdxi4525m ^ cdxi1799m);
wire cdxi4527m = reg_0_0&cdxi4526m;
wire cdxi4528m = a0&cdxi1597m;
wire cdxi4529m = reg_0_0&cdxi1614m;
wire cdxi4530m = a0&cdxi1701m;
wire cdxi4531m = reg_0_0&cdxi1718m;
wire cdxi4532m = cdxi2804m ^ r100m;
wire cdxi4533m = cdxi822m&cdxi208m;
wire cdxi4534m = cdxi362m&cdxi564m;
wire cdxi4535m = cdxi363m&cdxi778m;
wire cdxi4536m = cdxi825m&cdxi325m;
wire cdxi4537m = cdxi825m&cdxi326m;
wire cdxi4538m = cdxi1123m&r7m;
wire cdxi4539m = cdxi504m&cdxi430m;
wire cdxi4540m = cdxi938m&r9m;
wire cdxi4541m = cdxi822m&r12m;
wire cdxi4542m = cdxi1124m&r13m;
wire cdxi4543m = cdxi362m&cdxi567m;
wire cdxi4544m = cdxi362m&cdxi568m;
wire cdxi4545m = cdxi363m&cdxi781m;
wire cdxi4546m = cdxi363m&cdxi782m;
wire cdxi4547m = cdxi825m&r24m;
wire cdxi4548m = cdxi562m&r28m;
wire cdxi4549m = cdxi425m&r29m;
wire cdxi4550m = cdxi405m&r32m;
wire cdxi4551m = cdxi563m&r33m;
wire cdxi4552m = cdxi504m&r36m;
wire cdxi4553m = cdxi361m&r39m;
wire cdxi4554m = cdxi426m&r43m;
wire cdxi4555m = cdxi406m&r46m;
wire cdxi4556m = cdxi362m&r49m;
wire cdxi4557m = cdxi363m&r55m;
wire cdxi4558m = cdxi207m&r63m;
wire cdxi4559m = cdxi196m&r66m;
wire cdxi4560m = cdxi184m&r69m;
wire cdxi4561m = cdxi219m&r75m;
wire cdxi4562m = cdxi185m&r85m;
wire cdxi4563m = (cdxi4532m ^ cdxi4533m ^ cdxi4534m ^ cdxi4535m ^ cdxi4536m ^ cdxi4537m ^ cdxi4538m ^ cdxi4539m ^ cdxi4540m ^ cdxi4541m ^ cdxi4542m ^ cdxi4543m ^ cdxi4544m ^ cdxi4545m ^ cdxi4546m ^ cdxi4547m ^ cdxi4548m ^ cdxi4549m ^ cdxi4550m ^ cdxi4551m ^ cdxi4552m ^ cdxi4553m ^ cdxi4554m ^ cdxi4555m ^ cdxi4556m ^ cdxi4557m ^ cdxi4558m ^ cdxi4559m ^ cdxi4560m ^ cdxi4561m ^ cdxi4562m);
wire cdxi4564m = a0&cdxi4563m;
wire cdxi4565m = reg_0_2&cdxi1143m;
wire cdxi4566m = reg_0_1&cdxi1357m;
wire cdxi4567m = reg_0_1&cdxi1358m;
wire cdxi4568m = reg_0_1&cdxi1359m;
wire cdxi4569m = reg_0_1&cdxi1360m;
wire cdxi4570m = reg_0_3&cdxi3605m;
wire cdxi4571m = reg_0_2&cdxi1147m;
wire cdxi4572m = reg_0_2&cdxi1148m;
wire cdxi4573m = reg_0_2&cdxi1149m;
wire cdxi4574m = reg_0_1&cdxi1361m;
wire cdxi4575m = reg_0_1&cdxi1362m;
wire cdxi4576m = reg_0_1&cdxi1363m;
wire cdxi4577m = reg_0_1&cdxi1364m;
wire cdxi4578m = reg_0_1&cdxi1365m;
wire cdxi4579m = reg_0_1&cdxi1366m;
wire cdxi4580m = reg_0_4&cdxi970m;
wire cdxi4581m = reg_0_3&cdxi3611m;
wire cdxi4582m = reg_0_3&cdxi3612m;
wire cdxi4583m = reg_0_2&cdxi1153m;
wire cdxi4584m = reg_0_2&cdxi1154m;
wire cdxi4585m = reg_0_2&cdxi1155m;
wire cdxi4586m = reg_0_1&cdxi1367m;
wire cdxi4587m = reg_0_1&cdxi1368m;
wire cdxi4588m = reg_0_1&cdxi1369m;
wire cdxi4589m = reg_0_1&cdxi1370m;
wire cdxi4590m = reg_0_7&cdxi843m;
wire cdxi4591m = reg_0_4&cdxi959m;
wire cdxi4592m = reg_0_3&cdxi2150m;
wire cdxi4593m = reg_0_2&cdxi1142m;
wire cdxi4594m = reg_0_1&cdxi1356m;
wire cdxi4595m = (cdxi4565m ^ cdxi4566m ^ cdxi4567m ^ cdxi4568m ^ cdxi4569m ^ cdxi4570m ^ cdxi4571m ^ cdxi4572m ^ cdxi4573m ^ cdxi4574m ^ cdxi4575m ^ cdxi4576m ^ cdxi4577m ^ cdxi4578m ^ cdxi4579m ^ cdxi4580m ^ cdxi4581m ^ cdxi4582m ^ cdxi4583m ^ cdxi4584m ^ cdxi4585m ^ cdxi4586m ^ cdxi4587m ^ cdxi4588m ^ cdxi4589m ^ cdxi4590m ^ cdxi4591m ^ cdxi4592m ^ cdxi4593m ^ cdxi4594m ^ cdxi2871m);
wire cdxi4596m = reg_0_0&cdxi4595m;
wire cdxi4597m = 1&1 ^ cdxi184m ^ cdxi196m ^ cdxi240m ^ cdxi207m;
wire cdxi4598m = a0&cdxi4138m;
wire cdxi4599m = reg_0_0&cdxi4142m;
wire cdxi4600m = a0&cdxi293m;
wire cdxi4601m = reg_0_0&cdxi298m;
wire cdxi4602m = cdxi185m&cdxi253m;
wire cdxi4603m = reg_0_1&cdxi258m;
wire cdxi4604m = cdxi1763m ^ r67m;
wire cdxi4605m = cdxi219m&cdxi447m;
wire cdxi4606m = cdxi1233m&r1m;
wire cdxi4607m = cdxi363m&cdxi241m;
wire cdxi4608m = cdxi363m&cdxi242m;
wire cdxi4609m = cdxi445m&r7m;
wire cdxi4610m = cdxi219m&cdxi450m;
wire cdxi4611m = cdxi219m&cdxi451m;
wire cdxi4612m = cdxi446m&r14m;
wire cdxi4613m = cdxi406m&r15m;
wire cdxi4614m = cdxi363m&r22m;
wire cdxi4615m = cdxi240m&r29m;
wire cdxi4616m = cdxi196m&r30m;
wire cdxi4617m = cdxi219m&r37m;
wire cdxi4618m = cdxi185m&r47m;
wire cdxi4619m = (cdxi4604m ^ cdxi4605m ^ cdxi4606m ^ cdxi4607m ^ cdxi4608m ^ cdxi4609m ^ cdxi4610m ^ cdxi4611m ^ cdxi4612m ^ cdxi4613m ^ cdxi4614m ^ cdxi4615m ^ cdxi4616m ^ cdxi4617m ^ cdxi4618m);
wire cdxi4620m = a0&cdxi4619m;
wire cdxi4621m = reg_0_2&cdxi457m;
wire cdxi4622m = reg_0_1&cdxi535m;
wire cdxi4623m = reg_0_1&cdxi536m;
wire cdxi4624m = reg_0_1&cdxi537m;
wire cdxi4625m = reg_0_4&cdxi4457m;
wire cdxi4626m = reg_0_2&cdxi460m;
wire cdxi4627m = reg_0_2&cdxi461m;
wire cdxi4628m = reg_0_1&cdxi538m;
wire cdxi4629m = reg_0_1&cdxi539m;
wire cdxi4630m = reg_0_1&cdxi540m;
wire cdxi4631m = reg_0_5&cdxi842m;
wire cdxi4632m = reg_0_4&cdxi880m;
wire cdxi4633m = reg_0_2&cdxi456m;
wire cdxi4634m = reg_0_1&cdxi534m;
wire cdxi4635m = (cdxi4621m ^ cdxi4622m ^ cdxi4623m ^ cdxi4624m ^ cdxi4625m ^ cdxi4626m ^ cdxi4627m ^ cdxi4628m ^ cdxi4629m ^ cdxi4630m ^ cdxi4631m ^ cdxi4632m ^ cdxi4633m ^ cdxi4634m ^ cdxi1798m);
wire cdxi4636m = reg_0_0&cdxi4635m;
wire cdxi4637m = cdxi185m&cdxi1459m;
wire cdxi4638m = reg_0_1&cdxi1476m;
wire cdxi4639m = cdxi4062m;
wire cdxi4640m = 1&1 ^ a0 ^ cdxi184m ^ cdxi196m ^ cdxi218m ^ cdxi207m;
wire cdxi4641m = cdxi385m ^ r11m;
wire cdxi4642m = cdxi218m&r0m;
wire cdxi4643m = cdxi185m&r5m;
wire cdxi4644m = (cdxi4641m ^ cdxi4642m ^ cdxi4643m);
wire cdxi4645m = a0&cdxi4644m;
wire cdxi4646m = reg_0_6&cdxi130m;
wire cdxi4647m = reg_0_1&cdxi160m;
wire cdxi4648m = (cdxi4646m ^ cdxi4647m ^ cdxi394m);
wire cdxi4649m = reg_0_0&cdxi4648m;
wire cdxi4650m = 1&1 ^ a0 ^ cdxi185m ^ cdxi196m ^ cdxi218m;
wire cdxi4651m = a0&cdxi764m;
wire cdxi4652m = reg_0_0&cdxi773m;
wire cdxi4653m = cdxi219m&cdxi645m;
wire cdxi4654m = reg_0_2&cdxi654m;
wire cdxi4655m = cdxi185m&cdxi1354m;
wire cdxi4656m = reg_0_1&cdxi1371m;
wire cdxi4657m = cdxi1124m ^ r39m;
wire cdxi4658m = cdxi1905m ^ r76m;
wire cdxi4659m = cdxi3078m ^ r105m;
wire cdxi4660m = cdxi2801m ^ r110m;
wire cdxi4661m = 0&0 ^ a1 ^ b1 ^ c1 ^ f1;
wire cdxi4662m = b1 ^ r0m;
wire cdxi4663m = a1&cdxi0m;
wire cdxi4664m = (reg_1_8);
wire cdxi4665m = (cdxi4664m);
wire cdxi4666m = reg_1_0&cdxi4665m;
wire cdxi4667m = c1 ^ r1m;
wire cdxi4668m = a1&cdxi1m;
wire cdxi4669m = (reg_1_9);
wire cdxi4670m = (cdxi4669m);
wire cdxi4671m = reg_1_0&cdxi4670m;
wire cdxi4672m = d1 ^ r2m;
wire cdxi4673m = a1&cdxi2m;
wire cdxi4674m = (reg_1_10);
wire cdxi4675m = (cdxi4674m);
wire cdxi4676m = reg_1_0&cdxi4675m;
wire cdxi4677m = e1 ^ r3m;
wire cdxi4678m = a1&cdxi3m;
wire cdxi4679m = (reg_1_11);
wire cdxi4680m = (cdxi4679m);
wire cdxi4681m = reg_1_0&cdxi4680m;
wire cdxi4682m = f1 ^ r4m;
wire cdxi4683m = a1&cdxi4m;
wire cdxi4684m = (reg_1_12);
wire cdxi4685m = (cdxi4684m);
wire cdxi4686m = reg_1_0&cdxi4685m;
wire cdxi4687m = g1 ^ r5m;
wire cdxi4688m = a1&cdxi5m;
wire cdxi4689m = (reg_1_13);
wire cdxi4690m = (cdxi4689m);
wire cdxi4691m = reg_1_0&cdxi4690m;
wire cdxi4692m = b1&cdxi2m;
wire cdxi4693m = reg_1_1&cdxi4675m;
wire cdxi4694m = b1&cdxi5m;
wire cdxi4695m = reg_1_1&cdxi4690m;
wire cdxi4696m = h1 ^ r6m;
wire cdxi4697m = b1&cdxi6m;
wire cdxi4698m = (reg_1_14);
wire cdxi4699m = (cdxi4698m);
wire cdxi4700m = reg_1_1&cdxi4699m;
wire cdxi4701m = c1&cdxi5m;
wire cdxi4702m = reg_1_2&cdxi4690m;
wire cdxi4703m = d1&cdxi4m;
wire cdxi4704m = reg_1_3&cdxi4685m;
wire cdxi4705m = e1&cdxi5m;
wire cdxi4706m = reg_1_4&cdxi4690m;
wire cdxi4707m = e1&cdxi6m;
wire cdxi4708m = reg_1_4&cdxi4699m;
wire cdxi4709m = f1&cdxi5m;
wire cdxi4710m = reg_1_5&cdxi4690m;
wire cdxi4711m = d1;
wire cdxi4712m = b1;
wire cdxi4713m = cdxi4711m&r0m;
wire cdxi4714m = cdxi4712m&r2m;
wire cdxi4715m = (cdxi8m ^ cdxi4713m ^ cdxi4714m);
wire cdxi4716m = a1&cdxi4715m;
wire cdxi4717m = (reg_1_16);
wire cdxi4718m = reg_1_3&cdxi4664m;
wire cdxi4719m = reg_1_1&cdxi4674m;
wire cdxi4720m = (cdxi4718m ^ cdxi4719m ^ cdxi4717m);
wire cdxi4721m = reg_1_0&cdxi4720m;
wire cdxi4722m = e1;
wire cdxi4723m = cdxi4722m&r0m;
wire cdxi4724m = cdxi4712m&r3m;
wire cdxi4725m = (cdxi9m ^ cdxi4723m ^ cdxi4724m);
wire cdxi4726m = a1&cdxi4725m;
wire cdxi4727m = (reg_1_17);
wire cdxi4728m = reg_1_4&cdxi4664m;
wire cdxi4729m = reg_1_1&cdxi4679m;
wire cdxi4730m = (cdxi4728m ^ cdxi4729m ^ cdxi4727m);
wire cdxi4731m = reg_1_0&cdxi4730m;
wire cdxi4732m = h1;
wire cdxi4733m = cdxi4732m&r0m;
wire cdxi4734m = cdxi4712m&r6m;
wire cdxi4735m = (cdxi12m ^ cdxi4733m ^ cdxi4734m);
wire cdxi4736m = a1&cdxi4735m;
wire cdxi4737m = (reg_1_20);
wire cdxi4738m = reg_1_7&cdxi4664m;
wire cdxi4739m = reg_1_1&cdxi4698m;
wire cdxi4740m = (cdxi4738m ^ cdxi4739m ^ cdxi4737m);
wire cdxi4741m = reg_1_0&cdxi4740m;
wire cdxi4742m = g1;
wire cdxi4743m = c1;
wire cdxi4744m = cdxi4742m&r1m;
wire cdxi4745m = cdxi4743m&r5m;
wire cdxi4746m = (cdxi16m ^ cdxi4744m ^ cdxi4745m);
wire cdxi4747m = a1&cdxi4746m;
wire cdxi4748m = (reg_1_24);
wire cdxi4749m = reg_1_6&cdxi4669m;
wire cdxi4750m = reg_1_2&cdxi4689m;
wire cdxi4751m = (cdxi4749m ^ cdxi4750m ^ cdxi4748m);
wire cdxi4752m = reg_1_0&cdxi4751m;
wire cdxi4753m = cdxi4732m&r2m;
wire cdxi4754m = cdxi4711m&r6m;
wire cdxi4755m = (cdxi21m ^ cdxi4753m ^ cdxi4754m);
wire cdxi4756m = a1&cdxi4755m;
wire cdxi4757m = (reg_1_29);
wire cdxi4758m = reg_1_7&cdxi4674m;
wire cdxi4759m = reg_1_3&cdxi4698m;
wire cdxi4760m = (cdxi4758m ^ cdxi4759m ^ cdxi4757m);
wire cdxi4761m = reg_1_0&cdxi4760m;
wire cdxi4762m = f1;
wire cdxi4763m = cdxi4762m&r3m;
wire cdxi4764m = cdxi4722m&r4m;
wire cdxi4765m = (cdxi22m ^ cdxi4763m ^ cdxi4764m);
wire cdxi4766m = a1&cdxi4765m;
wire cdxi4767m = (reg_1_30);
wire cdxi4768m = reg_1_5&cdxi4679m;
wire cdxi4769m = reg_1_4&cdxi4684m;
wire cdxi4770m = (cdxi4768m ^ cdxi4769m ^ cdxi4767m);
wire cdxi4771m = reg_1_0&cdxi4770m;
wire cdxi4772m = cdxi4742m&r4m;
wire cdxi4773m = cdxi4762m&r5m;
wire cdxi4774m = (cdxi25m ^ cdxi4772m ^ cdxi4773m);
wire cdxi4775m = a1&cdxi4774m;
wire cdxi4776m = (reg_1_33);
wire cdxi4777m = reg_1_6&cdxi4684m;
wire cdxi4778m = reg_1_5&cdxi4689m;
wire cdxi4779m = (cdxi4777m ^ cdxi4778m ^ cdxi4776m);
wire cdxi4780m = reg_1_0&cdxi4779m;
wire cdxi4781m = cdxi4732m&r4m;
wire cdxi4782m = cdxi4762m&r6m;
wire cdxi4783m = (cdxi26m ^ cdxi4781m ^ cdxi4782m);
wire cdxi4784m = a1&cdxi4783m;
wire cdxi4785m = (reg_1_34);
wire cdxi4786m = reg_1_7&cdxi4684m;
wire cdxi4787m = reg_1_5&cdxi4698m;
wire cdxi4788m = (cdxi4786m ^ cdxi4787m ^ cdxi4785m);
wire cdxi4789m = reg_1_0&cdxi4788m;
wire cdxi4790m = cdxi4732m&r1m;
wire cdxi4791m = cdxi4743m&r6m;
wire cdxi4792m = (cdxi17m ^ cdxi4790m ^ cdxi4791m);
wire cdxi4793m = cdxi4712m&cdxi4792m;
wire cdxi4794m = (reg_1_25);
wire cdxi4795m = reg_1_7&cdxi4669m;
wire cdxi4796m = reg_1_2&cdxi4698m;
wire cdxi4797m = (cdxi4795m ^ cdxi4796m ^ cdxi4794m);
wire cdxi4798m = reg_1_1&cdxi4797m;
wire cdxi4799m = cdxi4722m&r2m;
wire cdxi4800m = cdxi4711m&r3m;
wire cdxi4801m = (cdxi18m ^ cdxi4799m ^ cdxi4800m);
wire cdxi4802m = cdxi4712m&cdxi4801m;
wire cdxi4803m = (reg_1_26);
wire cdxi4804m = reg_1_4&cdxi4674m;
wire cdxi4805m = reg_1_3&cdxi4679m;
wire cdxi4806m = (cdxi4804m ^ cdxi4805m ^ cdxi4803m);
wire cdxi4807m = reg_1_1&cdxi4806m;
wire cdxi4808m = cdxi4742m&r2m;
wire cdxi4809m = cdxi4711m&r5m;
wire cdxi4810m = (cdxi20m ^ cdxi4808m ^ cdxi4809m);
wire cdxi4811m = cdxi4712m&cdxi4810m;
wire cdxi4812m = (reg_1_28);
wire cdxi4813m = reg_1_6&cdxi4674m;
wire cdxi4814m = reg_1_3&cdxi4689m;
wire cdxi4815m = (cdxi4813m ^ cdxi4814m ^ cdxi4812m);
wire cdxi4816m = reg_1_1&cdxi4815m;
wire cdxi4817m = cdxi4742m&r3m;
wire cdxi4818m = cdxi4722m&r5m;
wire cdxi4819m = (cdxi23m ^ cdxi4817m ^ cdxi4818m);
wire cdxi4820m = cdxi4712m&cdxi4819m;
wire cdxi4821m = (reg_1_31);
wire cdxi4822m = reg_1_6&cdxi4679m;
wire cdxi4823m = reg_1_4&cdxi4689m;
wire cdxi4824m = (cdxi4822m ^ cdxi4823m ^ cdxi4821m);
wire cdxi4825m = reg_1_1&cdxi4824m;
wire cdxi4826m = cdxi4762m&r2m;
wire cdxi4827m = cdxi4711m&r4m;
wire cdxi4828m = (cdxi19m ^ cdxi4826m ^ cdxi4827m);
wire cdxi4829m = cdxi4743m&cdxi4828m;
wire cdxi4830m = (reg_1_27);
wire cdxi4831m = reg_1_5&cdxi4674m;
wire cdxi4832m = reg_1_3&cdxi4684m;
wire cdxi4833m = (cdxi4831m ^ cdxi4832m ^ cdxi4830m);
wire cdxi4834m = reg_1_2&cdxi4833m;
wire cdxi4835m = cdxi4743m&cdxi4755m;
wire cdxi4836m = reg_1_2&cdxi4760m;
wire cdxi4837m = cdxi4743m&cdxi4819m;
wire cdxi4838m = reg_1_2&cdxi4824m;
wire cdxi4839m = cdxi4732m&r3m;
wire cdxi4840m = cdxi4722m&r6m;
wire cdxi4841m = (cdxi24m ^ cdxi4839m ^ cdxi4840m);
wire cdxi4842m = cdxi4743m&cdxi4841m;
wire cdxi4843m = (reg_1_32);
wire cdxi4844m = reg_1_7&cdxi4679m;
wire cdxi4845m = reg_1_4&cdxi4698m;
wire cdxi4846m = (cdxi4844m ^ cdxi4845m ^ cdxi4843m);
wire cdxi4847m = reg_1_2&cdxi4846m;
wire cdxi4848m = cdxi4743m&cdxi4774m;
wire cdxi4849m = reg_1_2&cdxi4779m;
wire cdxi4850m = cdxi4732m&r5m;
wire cdxi4851m = cdxi4742m&r6m;
wire cdxi4852m = (cdxi27m ^ cdxi4850m ^ cdxi4851m);
wire cdxi4853m = cdxi4743m&cdxi4852m;
wire cdxi4854m = (reg_1_35);
wire cdxi4855m = reg_1_7&cdxi4689m;
wire cdxi4856m = reg_1_6&cdxi4698m;
wire cdxi4857m = (cdxi4855m ^ cdxi4856m ^ cdxi4854m);
wire cdxi4858m = reg_1_2&cdxi4857m;
wire cdxi4859m = cdxi4711m&cdxi4765m;
wire cdxi4860m = reg_1_3&cdxi4770m;
wire cdxi4861m = cdxi4711m&cdxi4819m;
wire cdxi4862m = reg_1_3&cdxi4824m;
wire cdxi4863m = cdxi4711m&cdxi4841m;
wire cdxi4864m = reg_1_3&cdxi4846m;
wire cdxi4865m = cdxi4711m&cdxi4774m;
wire cdxi4866m = reg_1_3&cdxi4779m;
wire cdxi4867m = cdxi4711m&cdxi4783m;
wire cdxi4868m = reg_1_3&cdxi4788m;
wire cdxi4869m = cdxi4722m&cdxi4774m;
wire cdxi4870m = reg_1_4&cdxi4779m;
wire cdxi4871m = cdxi4722m&cdxi4783m;
wire cdxi4872m = reg_1_4&cdxi4788m;
wire cdxi4873m = cdxi4743m&cdxi4711m;
wire cdxi4874m = cdxi4712m&cdxi4711m;
wire cdxi4875m = cdxi4712m&cdxi4743m;
wire cdxi4876m = cdxi4743m&cdxi4713m;
wire cdxi4877m = cdxi4874m&r1m;
wire cdxi4878m = cdxi4875m&r2m;
wire cdxi4879m = cdxi4711m&r7m;
wire cdxi4880m = cdxi4743m&r8m;
wire cdxi4881m = cdxi4712m&r13m;
wire cdxi4882m = (cdxi28m ^ cdxi4876m ^ cdxi4877m ^ cdxi4878m ^ cdxi4879m ^ cdxi4880m ^ cdxi4881m);
wire cdxi4883m = a1&cdxi4882m;
wire cdxi4884m = (reg_1_15);
wire cdxi4885m = (reg_1_21);
wire cdxi4886m = (reg_1_36);
wire cdxi4887m = reg_1_2&cdxi4718m;
wire cdxi4888m = reg_1_1&reg_1_3&cdxi4669m;
wire cdxi4889m = reg_1_1&reg_1_2&cdxi4674m;
wire cdxi4890m = reg_1_3&cdxi4884m;
wire cdxi4891m = reg_1_2&cdxi4717m;
wire cdxi4892m = reg_1_1&cdxi4885m;
wire cdxi4893m = (cdxi4887m ^ cdxi4888m ^ cdxi4889m ^ cdxi4890m ^ cdxi4891m ^ cdxi4892m ^ cdxi4886m);
wire cdxi4894m = reg_1_0&cdxi4893m;
wire cdxi4895m = cdxi4743m&cdxi4742m;
wire cdxi4896m = cdxi4712m&cdxi4742m;
wire cdxi4897m = cdxi4895m&r0m;
wire cdxi4898m = cdxi4712m&cdxi4744m;
wire cdxi4899m = cdxi4712m&cdxi4745m;
wire cdxi4900m = cdxi4742m&r7m;
wire cdxi4901m = cdxi4743m&r11m;
wire cdxi4902m = cdxi4712m&r16m;
wire cdxi4903m = (cdxi31m ^ cdxi4897m ^ cdxi4898m ^ cdxi4899m ^ cdxi4900m ^ cdxi4901m ^ cdxi4902m);
wire cdxi4904m = a1&cdxi4903m;
wire cdxi4905m = (reg_1_19);
wire cdxi4906m = (reg_1_39);
wire cdxi4907m = reg_1_2&reg_1_6&cdxi4664m;
wire cdxi4908m = reg_1_1&cdxi4749m;
wire cdxi4909m = reg_1_1&cdxi4750m;
wire cdxi4910m = reg_1_6&cdxi4884m;
wire cdxi4911m = reg_1_2&cdxi4905m;
wire cdxi4912m = reg_1_1&cdxi4748m;
wire cdxi4913m = (cdxi4907m ^ cdxi4908m ^ cdxi4909m ^ cdxi4910m ^ cdxi4911m ^ cdxi4912m ^ cdxi4906m);
wire cdxi4914m = reg_1_0&cdxi4913m;
wire cdxi4915m = cdxi4711m&cdxi4722m;
wire cdxi4916m = cdxi4712m&cdxi4722m;
wire cdxi4917m = cdxi4711m&cdxi4723m;
wire cdxi4918m = cdxi4712m&cdxi4799m;
wire cdxi4919m = cdxi4712m&cdxi4800m;
wire cdxi4920m = cdxi4722m&r8m;
wire cdxi4921m = cdxi4711m&r9m;
wire cdxi4922m = cdxi4712m&r18m;
wire cdxi4923m = (cdxi33m ^ cdxi4917m ^ cdxi4918m ^ cdxi4919m ^ cdxi4920m ^ cdxi4921m ^ cdxi4922m);
wire cdxi4924m = a1&cdxi4923m;
wire cdxi4925m = (reg_1_41);
wire cdxi4926m = reg_1_3&cdxi4728m;
wire cdxi4927m = reg_1_1&cdxi4804m;
wire cdxi4928m = reg_1_1&cdxi4805m;
wire cdxi4929m = reg_1_4&cdxi4717m;
wire cdxi4930m = reg_1_3&cdxi4727m;
wire cdxi4931m = reg_1_1&cdxi4803m;
wire cdxi4932m = (cdxi4926m ^ cdxi4927m ^ cdxi4928m ^ cdxi4929m ^ cdxi4930m ^ cdxi4931m ^ cdxi4925m);
wire cdxi4933m = reg_1_0&cdxi4932m;
wire cdxi4934m = cdxi4711m&cdxi4732m;
wire cdxi4935m = cdxi4712m&cdxi4732m;
wire cdxi4936m = cdxi4711m&cdxi4733m;
wire cdxi4937m = cdxi4712m&cdxi4753m;
wire cdxi4938m = cdxi4712m&cdxi4754m;
wire cdxi4939m = cdxi4732m&r8m;
wire cdxi4940m = cdxi4711m&r12m;
wire cdxi4941m = cdxi4712m&r21m;
wire cdxi4942m = (cdxi36m ^ cdxi4936m ^ cdxi4937m ^ cdxi4938m ^ cdxi4939m ^ cdxi4940m ^ cdxi4941m);
wire cdxi4943m = a1&cdxi4942m;
wire cdxi4944m = (reg_1_44);
wire cdxi4945m = reg_1_3&cdxi4738m;
wire cdxi4946m = reg_1_1&cdxi4758m;
wire cdxi4947m = reg_1_1&cdxi4759m;
wire cdxi4948m = reg_1_7&cdxi4717m;
wire cdxi4949m = reg_1_3&cdxi4737m;
wire cdxi4950m = reg_1_1&cdxi4757m;
wire cdxi4951m = (cdxi4945m ^ cdxi4946m ^ cdxi4947m ^ cdxi4948m ^ cdxi4949m ^ cdxi4950m ^ cdxi4944m);
wire cdxi4952m = reg_1_0&cdxi4951m;
wire cdxi4953m = cdxi4722m&cdxi4762m;
wire cdxi4954m = cdxi4712m&cdxi4762m;
wire cdxi4955m = cdxi4953m&r0m;
wire cdxi4956m = cdxi4712m&cdxi4763m;
wire cdxi4957m = cdxi4712m&cdxi4764m;
wire cdxi4958m = cdxi4762m&r9m;
wire cdxi4959m = cdxi4722m&r10m;
wire cdxi4960m = cdxi4712m&r22m;
wire cdxi4961m = (cdxi37m ^ cdxi4955m ^ cdxi4956m ^ cdxi4957m ^ cdxi4958m ^ cdxi4959m ^ cdxi4960m);
wire cdxi4962m = a1&cdxi4961m;
wire cdxi4963m = (reg_1_18);
wire cdxi4964m = (reg_1_45);
wire cdxi4965m = reg_1_4&reg_1_5&cdxi4664m;
wire cdxi4966m = reg_1_1&cdxi4768m;
wire cdxi4967m = reg_1_1&cdxi4769m;
wire cdxi4968m = reg_1_5&cdxi4727m;
wire cdxi4969m = reg_1_4&cdxi4963m;
wire cdxi4970m = reg_1_1&cdxi4767m;
wire cdxi4971m = (cdxi4965m ^ cdxi4966m ^ cdxi4967m ^ cdxi4968m ^ cdxi4969m ^ cdxi4970m ^ cdxi4964m);
wire cdxi4972m = reg_1_0&cdxi4971m;
wire cdxi4973m = cdxi4722m&cdxi4742m;
wire cdxi4974m = cdxi4973m&r0m;
wire cdxi4975m = cdxi4712m&cdxi4817m;
wire cdxi4976m = cdxi4712m&cdxi4818m;
wire cdxi4977m = cdxi4742m&r9m;
wire cdxi4978m = cdxi4722m&r11m;
wire cdxi4979m = cdxi4712m&r23m;
wire cdxi4980m = (cdxi38m ^ cdxi4974m ^ cdxi4975m ^ cdxi4976m ^ cdxi4977m ^ cdxi4978m ^ cdxi4979m);
wire cdxi4981m = a1&cdxi4980m;
wire cdxi4982m = (reg_1_46);
wire cdxi4983m = reg_1_4&reg_1_6&cdxi4664m;
wire cdxi4984m = reg_1_1&cdxi4822m;
wire cdxi4985m = reg_1_1&cdxi4823m;
wire cdxi4986m = reg_1_6&cdxi4727m;
wire cdxi4987m = reg_1_4&cdxi4905m;
wire cdxi4988m = reg_1_1&cdxi4821m;
wire cdxi4989m = (cdxi4983m ^ cdxi4984m ^ cdxi4985m ^ cdxi4986m ^ cdxi4987m ^ cdxi4988m ^ cdxi4982m);
wire cdxi4990m = reg_1_0&cdxi4989m;
wire cdxi4991m = cdxi4762m&cdxi4732m;
wire cdxi4992m = cdxi4762m&cdxi4733m;
wire cdxi4993m = cdxi4712m&cdxi4781m;
wire cdxi4994m = cdxi4712m&cdxi4782m;
wire cdxi4995m = cdxi4732m&r10m;
wire cdxi4996m = cdxi4762m&r12m;
wire cdxi4997m = cdxi4712m&r26m;
wire cdxi4998m = (cdxi41m ^ cdxi4992m ^ cdxi4993m ^ cdxi4994m ^ cdxi4995m ^ cdxi4996m ^ cdxi4997m);
wire cdxi4999m = a1&cdxi4998m;
wire cdxi5000m = (reg_1_49);
wire cdxi5001m = reg_1_5&cdxi4738m;
wire cdxi5002m = reg_1_1&cdxi4786m;
wire cdxi5003m = reg_1_1&cdxi4787m;
wire cdxi5004m = reg_1_7&cdxi4963m;
wire cdxi5005m = reg_1_5&cdxi4737m;
wire cdxi5006m = reg_1_1&cdxi4785m;
wire cdxi5007m = (cdxi5001m ^ cdxi5002m ^ cdxi5003m ^ cdxi5004m ^ cdxi5005m ^ cdxi5006m ^ cdxi5000m);
wire cdxi5008m = reg_1_0&cdxi5007m;
wire cdxi5009m = cdxi4743m&cdxi4722m;
wire cdxi5010m = cdxi4915m&r1m;
wire cdxi5011m = cdxi4743m&cdxi4799m;
wire cdxi5012m = cdxi4743m&cdxi4800m;
wire cdxi5013m = cdxi4722m&r13m;
wire cdxi5014m = cdxi4711m&r14m;
wire cdxi5015m = cdxi4743m&r18m;
wire cdxi5016m = (cdxi43m ^ cdxi5010m ^ cdxi5011m ^ cdxi5012m ^ cdxi5013m ^ cdxi5014m ^ cdxi5015m);
wire cdxi5017m = a1&cdxi5016m;
wire cdxi5018m = (reg_1_22);
wire cdxi5019m = (reg_1_51);
wire cdxi5020m = reg_1_3&reg_1_4&cdxi4669m;
wire cdxi5021m = reg_1_2&cdxi4804m;
wire cdxi5022m = reg_1_2&cdxi4805m;
wire cdxi5023m = reg_1_4&cdxi4885m;
wire cdxi5024m = reg_1_3&cdxi5018m;
wire cdxi5025m = reg_1_2&cdxi4803m;
wire cdxi5026m = (cdxi5020m ^ cdxi5021m ^ cdxi5022m ^ cdxi5023m ^ cdxi5024m ^ cdxi5025m ^ cdxi5019m);
wire cdxi5027m = reg_1_0&cdxi5026m;
wire cdxi5028m = cdxi4743m&cdxi4762m;
wire cdxi5029m = cdxi4953m&r1m;
wire cdxi5030m = cdxi4743m&cdxi4763m;
wire cdxi5031m = cdxi4743m&cdxi4764m;
wire cdxi5032m = cdxi4762m&r14m;
wire cdxi5033m = cdxi4722m&r15m;
wire cdxi5034m = cdxi4743m&r22m;
wire cdxi5035m = (cdxi47m ^ cdxi5029m ^ cdxi5030m ^ cdxi5031m ^ cdxi5032m ^ cdxi5033m ^ cdxi5034m);
wire cdxi5036m = a1&cdxi5035m;
wire cdxi5037m = (reg_1_23);
wire cdxi5038m = (reg_1_55);
wire cdxi5039m = reg_1_4&reg_1_5&cdxi4669m;
wire cdxi5040m = reg_1_2&cdxi4768m;
wire cdxi5041m = reg_1_2&cdxi4769m;
wire cdxi5042m = reg_1_5&cdxi5018m;
wire cdxi5043m = reg_1_4&cdxi5037m;
wire cdxi5044m = reg_1_2&cdxi4767m;
wire cdxi5045m = (cdxi5039m ^ cdxi5040m ^ cdxi5041m ^ cdxi5042m ^ cdxi5043m ^ cdxi5044m ^ cdxi5038m);
wire cdxi5046m = reg_1_0&cdxi5045m;
wire cdxi5047m = cdxi4722m&cdxi4744m;
wire cdxi5048m = cdxi4743m&cdxi4817m;
wire cdxi5049m = cdxi4743m&cdxi4818m;
wire cdxi5050m = cdxi4742m&r14m;
wire cdxi5051m = cdxi4722m&r16m;
wire cdxi5052m = cdxi4743m&r23m;
wire cdxi5053m = (cdxi48m ^ cdxi5047m ^ cdxi5048m ^ cdxi5049m ^ cdxi5050m ^ cdxi5051m ^ cdxi5052m);
wire cdxi5054m = a1&cdxi5053m;
wire cdxi5055m = (reg_1_56);
wire cdxi5056m = reg_1_4&cdxi4749m;
wire cdxi5057m = reg_1_2&cdxi4822m;
wire cdxi5058m = reg_1_2&cdxi4823m;
wire cdxi5059m = reg_1_6&cdxi5018m;
wire cdxi5060m = reg_1_4&cdxi4748m;
wire cdxi5061m = reg_1_2&cdxi4821m;
wire cdxi5062m = (cdxi5056m ^ cdxi5057m ^ cdxi5058m ^ cdxi5059m ^ cdxi5060m ^ cdxi5061m ^ cdxi5055m);
wire cdxi5063m = reg_1_0&cdxi5062m;
wire cdxi5064m = cdxi4722m&cdxi4732m;
wire cdxi5065m = cdxi4743m&cdxi4732m;
wire cdxi5066m = cdxi4722m&cdxi4790m;
wire cdxi5067m = cdxi4743m&cdxi4839m;
wire cdxi5068m = cdxi4743m&cdxi4840m;
wire cdxi5069m = cdxi4732m&r14m;
wire cdxi5070m = cdxi4722m&r17m;
wire cdxi5071m = cdxi4743m&r24m;
wire cdxi5072m = (cdxi49m ^ cdxi5066m ^ cdxi5067m ^ cdxi5068m ^ cdxi5069m ^ cdxi5070m ^ cdxi5071m);
wire cdxi5073m = a1&cdxi5072m;
wire cdxi5074m = (reg_1_57);
wire cdxi5075m = reg_1_4&cdxi4795m;
wire cdxi5076m = reg_1_2&cdxi4844m;
wire cdxi5077m = reg_1_2&cdxi4845m;
wire cdxi5078m = reg_1_7&cdxi5018m;
wire cdxi5079m = reg_1_4&cdxi4794m;
wire cdxi5080m = reg_1_2&cdxi4843m;
wire cdxi5081m = (cdxi5075m ^ cdxi5076m ^ cdxi5077m ^ cdxi5078m ^ cdxi5079m ^ cdxi5080m ^ cdxi5074m);
wire cdxi5082m = reg_1_0&cdxi5081m;
wire cdxi5083m = cdxi4711m&cdxi4762m;
wire cdxi5084m = cdxi4722m&cdxi4826m;
wire cdxi5085m = cdxi4711m&cdxi4763m;
wire cdxi5086m = cdxi4711m&cdxi4764m;
wire cdxi5087m = cdxi4762m&r18m;
wire cdxi5088m = cdxi4722m&r19m;
wire cdxi5089m = cdxi4711m&r22m;
wire cdxi5090m = (cdxi53m ^ cdxi5084m ^ cdxi5085m ^ cdxi5086m ^ cdxi5087m ^ cdxi5088m ^ cdxi5089m);
wire cdxi5091m = a1&cdxi5090m;
wire cdxi5092m = (reg_1_61);
wire cdxi5093m = reg_1_4&cdxi4831m;
wire cdxi5094m = reg_1_3&cdxi4768m;
wire cdxi5095m = reg_1_3&cdxi4769m;
wire cdxi5096m = reg_1_5&cdxi4803m;
wire cdxi5097m = reg_1_4&cdxi4830m;
wire cdxi5098m = reg_1_3&cdxi4767m;
wire cdxi5099m = (cdxi5093m ^ cdxi5094m ^ cdxi5095m ^ cdxi5096m ^ cdxi5097m ^ cdxi5098m ^ cdxi5092m);
wire cdxi5100m = reg_1_0&cdxi5099m;
wire cdxi5101m = cdxi4711m&cdxi4742m;
wire cdxi5102m = cdxi4722m&cdxi4808m;
wire cdxi5103m = cdxi4711m&cdxi4817m;
wire cdxi5104m = cdxi4711m&cdxi4818m;
wire cdxi5105m = cdxi4742m&r18m;
wire cdxi5106m = cdxi4722m&r20m;
wire cdxi5107m = cdxi4711m&r23m;
wire cdxi5108m = (cdxi54m ^ cdxi5102m ^ cdxi5103m ^ cdxi5104m ^ cdxi5105m ^ cdxi5106m ^ cdxi5107m);
wire cdxi5109m = a1&cdxi5108m;
wire cdxi5110m = (reg_1_62);
wire cdxi5111m = reg_1_4&cdxi4813m;
wire cdxi5112m = reg_1_3&cdxi4822m;
wire cdxi5113m = reg_1_3&cdxi4823m;
wire cdxi5114m = reg_1_6&cdxi4803m;
wire cdxi5115m = reg_1_4&cdxi4812m;
wire cdxi5116m = reg_1_3&cdxi4821m;
wire cdxi5117m = (cdxi5111m ^ cdxi5112m ^ cdxi5113m ^ cdxi5114m ^ cdxi5115m ^ cdxi5116m ^ cdxi5110m);
wire cdxi5118m = reg_1_0&cdxi5117m;
wire cdxi5119m = cdxi4762m&cdxi4753m;
wire cdxi5120m = cdxi4711m&cdxi4781m;
wire cdxi5121m = cdxi4711m&cdxi4782m;
wire cdxi5122m = cdxi4732m&r19m;
wire cdxi5123m = cdxi4762m&r21m;
wire cdxi5124m = cdxi4711m&r26m;
wire cdxi5125m = (cdxi57m ^ cdxi5119m ^ cdxi5120m ^ cdxi5121m ^ cdxi5122m ^ cdxi5123m ^ cdxi5124m);
wire cdxi5126m = a1&cdxi5125m;
wire cdxi5127m = (reg_1_65);
wire cdxi5128m = reg_1_5&cdxi4758m;
wire cdxi5129m = reg_1_3&cdxi4786m;
wire cdxi5130m = reg_1_3&cdxi4787m;
wire cdxi5131m = reg_1_7&cdxi4830m;
wire cdxi5132m = reg_1_5&cdxi4757m;
wire cdxi5133m = reg_1_3&cdxi4785m;
wire cdxi5134m = (cdxi5128m ^ cdxi5129m ^ cdxi5130m ^ cdxi5131m ^ cdxi5132m ^ cdxi5133m ^ cdxi5127m);
wire cdxi5135m = reg_1_0&cdxi5134m;
wire cdxi5136m = cdxi4762m&cdxi4742m;
wire cdxi5137m = cdxi4762m&cdxi4817m;
wire cdxi5138m = cdxi4722m&cdxi4772m;
wire cdxi5139m = cdxi4722m&cdxi4773m;
wire cdxi5140m = cdxi4742m&r22m;
wire cdxi5141m = cdxi4762m&r23m;
wire cdxi5142m = cdxi4722m&r25m;
wire cdxi5143m = (cdxi59m ^ cdxi5137m ^ cdxi5138m ^ cdxi5139m ^ cdxi5140m ^ cdxi5141m ^ cdxi5142m);
wire cdxi5144m = a1&cdxi5143m;
wire cdxi5145m = (reg_1_67);
wire cdxi5146m = reg_1_5&cdxi4822m;
wire cdxi5147m = reg_1_4&cdxi4777m;
wire cdxi5148m = reg_1_4&cdxi4778m;
wire cdxi5149m = reg_1_6&cdxi4767m;
wire cdxi5150m = reg_1_5&cdxi4821m;
wire cdxi5151m = reg_1_4&cdxi4776m;
wire cdxi5152m = (cdxi5146m ^ cdxi5147m ^ cdxi5148m ^ cdxi5149m ^ cdxi5150m ^ cdxi5151m ^ cdxi5145m);
wire cdxi5153m = reg_1_0&cdxi5152m;
wire cdxi5154m = cdxi4742m&cdxi4732m;
wire cdxi5155m = cdxi4742m&cdxi4781m;
wire cdxi5156m = cdxi4762m&cdxi4850m;
wire cdxi5157m = cdxi4762m&cdxi4851m;
wire cdxi5158m = cdxi4732m&r25m;
wire cdxi5159m = cdxi4742m&r26m;
wire cdxi5160m = cdxi4762m&r27m;
wire cdxi5161m = (cdxi62m ^ cdxi5155m ^ cdxi5156m ^ cdxi5157m ^ cdxi5158m ^ cdxi5159m ^ cdxi5160m);
wire cdxi5162m = a1&cdxi5161m;
wire cdxi5163m = (reg_1_70);
wire cdxi5164m = reg_1_6&cdxi4786m;
wire cdxi5165m = reg_1_5&cdxi4855m;
wire cdxi5166m = reg_1_5&cdxi4856m;
wire cdxi5167m = reg_1_7&cdxi4776m;
wire cdxi5168m = reg_1_6&cdxi4785m;
wire cdxi5169m = reg_1_5&cdxi4854m;
wire cdxi5170m = (cdxi5164m ^ cdxi5165m ^ cdxi5166m ^ cdxi5167m ^ cdxi5168m ^ cdxi5169m ^ cdxi5163m);
wire cdxi5171m = reg_1_0&cdxi5170m;
wire cdxi5172m = cdxi5083m&r1m;
wire cdxi5173m = cdxi4743m&cdxi4826m;
wire cdxi5174m = cdxi4743m&cdxi4827m;
wire cdxi5175m = cdxi4762m&r13m;
wire cdxi5176m = cdxi4711m&r15m;
wire cdxi5177m = cdxi4743m&r19m;
wire cdxi5178m = (cdxi44m ^ cdxi5172m ^ cdxi5173m ^ cdxi5174m ^ cdxi5175m ^ cdxi5176m ^ cdxi5177m);
wire cdxi5179m = cdxi4712m&cdxi5178m;
wire cdxi5180m = (reg_1_52);
wire cdxi5181m = reg_1_3&reg_1_5&cdxi4669m;
wire cdxi5182m = reg_1_2&cdxi4831m;
wire cdxi5183m = reg_1_2&cdxi4832m;
wire cdxi5184m = reg_1_5&cdxi4885m;
wire cdxi5185m = reg_1_3&cdxi5037m;
wire cdxi5186m = reg_1_2&cdxi4830m;
wire cdxi5187m = (cdxi5181m ^ cdxi5182m ^ cdxi5183m ^ cdxi5184m ^ cdxi5185m ^ cdxi5186m ^ cdxi5180m);
wire cdxi5188m = reg_1_1&cdxi5187m;
wire cdxi5189m = cdxi4711m&cdxi4744m;
wire cdxi5190m = cdxi4743m&cdxi4808m;
wire cdxi5191m = cdxi4743m&cdxi4809m;
wire cdxi5192m = cdxi4742m&r13m;
wire cdxi5193m = cdxi4711m&r16m;
wire cdxi5194m = cdxi4743m&r20m;
wire cdxi5195m = (cdxi45m ^ cdxi5189m ^ cdxi5190m ^ cdxi5191m ^ cdxi5192m ^ cdxi5193m ^ cdxi5194m);
wire cdxi5196m = cdxi4712m&cdxi5195m;
wire cdxi5197m = (reg_1_53);
wire cdxi5198m = reg_1_3&cdxi4749m;
wire cdxi5199m = reg_1_2&cdxi4813m;
wire cdxi5200m = reg_1_2&cdxi4814m;
wire cdxi5201m = reg_1_6&cdxi4885m;
wire cdxi5202m = reg_1_3&cdxi4748m;
wire cdxi5203m = reg_1_2&cdxi4812m;
wire cdxi5204m = (cdxi5198m ^ cdxi5199m ^ cdxi5200m ^ cdxi5201m ^ cdxi5202m ^ cdxi5203m ^ cdxi5197m);
wire cdxi5205m = reg_1_1&cdxi5204m;
wire cdxi5206m = cdxi4712m&cdxi5053m;
wire cdxi5207m = reg_1_1&cdxi5062m;
wire cdxi5208m = cdxi4712m&cdxi5072m;
wire cdxi5209m = reg_1_1&cdxi5081m;
wire cdxi5210m = cdxi4762m&cdxi4744m;
wire cdxi5211m = cdxi4743m&cdxi4772m;
wire cdxi5212m = cdxi4743m&cdxi4773m;
wire cdxi5213m = cdxi4742m&r15m;
wire cdxi5214m = cdxi4762m&r16m;
wire cdxi5215m = cdxi4743m&r25m;
wire cdxi5216m = (cdxi50m ^ cdxi5210m ^ cdxi5211m ^ cdxi5212m ^ cdxi5213m ^ cdxi5214m ^ cdxi5215m);
wire cdxi5217m = cdxi4712m&cdxi5216m;
wire cdxi5218m = (reg_1_58);
wire cdxi5219m = reg_1_5&cdxi4749m;
wire cdxi5220m = reg_1_2&cdxi4777m;
wire cdxi5221m = reg_1_2&cdxi4778m;
wire cdxi5222m = reg_1_6&cdxi5037m;
wire cdxi5223m = reg_1_5&cdxi4748m;
wire cdxi5224m = reg_1_2&cdxi4776m;
wire cdxi5225m = (cdxi5219m ^ cdxi5220m ^ cdxi5221m ^ cdxi5222m ^ cdxi5223m ^ cdxi5224m ^ cdxi5218m);
wire cdxi5226m = reg_1_1&cdxi5225m;
wire cdxi5227m = cdxi4762m&cdxi4790m;
wire cdxi5228m = cdxi4743m&cdxi4781m;
wire cdxi5229m = cdxi4743m&cdxi4782m;
wire cdxi5230m = cdxi4732m&r15m;
wire cdxi5231m = cdxi4762m&r17m;
wire cdxi5232m = cdxi4743m&r26m;
wire cdxi5233m = (cdxi51m ^ cdxi5227m ^ cdxi5228m ^ cdxi5229m ^ cdxi5230m ^ cdxi5231m ^ cdxi5232m);
wire cdxi5234m = cdxi4712m&cdxi5233m;
wire cdxi5235m = (reg_1_59);
wire cdxi5236m = reg_1_5&cdxi4795m;
wire cdxi5237m = reg_1_2&cdxi4786m;
wire cdxi5238m = reg_1_2&cdxi4787m;
wire cdxi5239m = reg_1_7&cdxi5037m;
wire cdxi5240m = reg_1_5&cdxi4794m;
wire cdxi5241m = reg_1_2&cdxi4785m;
wire cdxi5242m = (cdxi5236m ^ cdxi5237m ^ cdxi5238m ^ cdxi5239m ^ cdxi5240m ^ cdxi5241m ^ cdxi5235m);
wire cdxi5243m = reg_1_1&cdxi5242m;
wire cdxi5244m = cdxi4712m&cdxi5090m;
wire cdxi5245m = reg_1_1&cdxi5099m;
wire cdxi5246m = cdxi4712m&cdxi5125m;
wire cdxi5247m = reg_1_1&cdxi5134m;
wire cdxi5248m = cdxi4712m&cdxi5143m;
wire cdxi5249m = reg_1_1&cdxi5152m;
wire cdxi5250m = cdxi4742m&cdxi4839m;
wire cdxi5251m = cdxi4722m&cdxi4850m;
wire cdxi5252m = cdxi4722m&cdxi4851m;
wire cdxi5253m = cdxi4732m&r23m;
wire cdxi5254m = cdxi4742m&r24m;
wire cdxi5255m = cdxi4722m&r27m;
wire cdxi5256m = (cdxi61m ^ cdxi5250m ^ cdxi5251m ^ cdxi5252m ^ cdxi5253m ^ cdxi5254m ^ cdxi5255m);
wire cdxi5257m = cdxi4712m&cdxi5256m;
wire cdxi5258m = (reg_1_69);
wire cdxi5259m = reg_1_6&cdxi4844m;
wire cdxi5260m = reg_1_4&cdxi4855m;
wire cdxi5261m = reg_1_4&cdxi4856m;
wire cdxi5262m = reg_1_7&cdxi4821m;
wire cdxi5263m = reg_1_6&cdxi4843m;
wire cdxi5264m = reg_1_4&cdxi4854m;
wire cdxi5265m = (cdxi5259m ^ cdxi5260m ^ cdxi5261m ^ cdxi5262m ^ cdxi5263m ^ cdxi5264m ^ cdxi5258m);
wire cdxi5266m = reg_1_1&cdxi5265m;
wire cdxi5267m = cdxi4743m&cdxi5090m;
wire cdxi5268m = reg_1_2&cdxi5099m;
wire cdxi5269m = cdxi4722m&cdxi4753m;
wire cdxi5270m = cdxi4711m&cdxi4839m;
wire cdxi5271m = cdxi4711m&cdxi4840m;
wire cdxi5272m = cdxi4732m&r18m;
wire cdxi5273m = cdxi4722m&r21m;
wire cdxi5274m = cdxi4711m&r24m;
wire cdxi5275m = (cdxi55m ^ cdxi5269m ^ cdxi5270m ^ cdxi5271m ^ cdxi5272m ^ cdxi5273m ^ cdxi5274m);
wire cdxi5276m = cdxi4743m&cdxi5275m;
wire cdxi5277m = (reg_1_63);
wire cdxi5278m = reg_1_4&cdxi4758m;
wire cdxi5279m = reg_1_3&cdxi4844m;
wire cdxi5280m = reg_1_3&cdxi4845m;
wire cdxi5281m = reg_1_7&cdxi4803m;
wire cdxi5282m = reg_1_4&cdxi4757m;
wire cdxi5283m = reg_1_3&cdxi4843m;
wire cdxi5284m = (cdxi5278m ^ cdxi5279m ^ cdxi5280m ^ cdxi5281m ^ cdxi5282m ^ cdxi5283m ^ cdxi5277m);
wire cdxi5285m = reg_1_2&cdxi5284m;
wire cdxi5286m = cdxi4743m&cdxi5125m;
wire cdxi5287m = reg_1_2&cdxi5134m;
wire cdxi5288m = cdxi4743m&cdxi5161m;
wire cdxi5289m = reg_1_2&cdxi5170m;
wire cdxi5290m = cdxi4711m&cdxi5143m;
wire cdxi5291m = reg_1_3&cdxi5152m;
wire cdxi5292m = cdxi4762m&cdxi4839m;
wire cdxi5293m = cdxi4722m&cdxi4781m;
wire cdxi5294m = cdxi4722m&cdxi4782m;
wire cdxi5295m = cdxi4732m&r22m;
wire cdxi5296m = cdxi4762m&r24m;
wire cdxi5297m = cdxi4722m&r26m;
wire cdxi5298m = (cdxi60m ^ cdxi5292m ^ cdxi5293m ^ cdxi5294m ^ cdxi5295m ^ cdxi5296m ^ cdxi5297m);
wire cdxi5299m = cdxi4711m&cdxi5298m;
wire cdxi5300m = (reg_1_68);
wire cdxi5301m = reg_1_5&cdxi4844m;
wire cdxi5302m = reg_1_4&cdxi4786m;
wire cdxi5303m = reg_1_4&cdxi4787m;
wire cdxi5304m = reg_1_7&cdxi4767m;
wire cdxi5305m = reg_1_5&cdxi4843m;
wire cdxi5306m = reg_1_4&cdxi4785m;
wire cdxi5307m = (cdxi5301m ^ cdxi5302m ^ cdxi5303m ^ cdxi5304m ^ cdxi5305m ^ cdxi5306m ^ cdxi5300m);
wire cdxi5308m = reg_1_3&cdxi5307m;
wire cdxi5309m = cdxi4711m&cdxi5256m;
wire cdxi5310m = reg_1_3&cdxi5265m;
wire cdxi5311m = cdxi4873m&cdxi4722m;
wire cdxi5312m = cdxi4874m&cdxi4722m;
wire cdxi5313m = cdxi4875m&cdxi4722m;
wire cdxi5314m = cdxi4712m&cdxi4873m;
wire cdxi5315m = cdxi4873m&cdxi4723m;
wire cdxi5316m = cdxi5312m&r1m;
wire cdxi5317m = cdxi4875m&cdxi4799m;
wire cdxi5318m = cdxi4875m&cdxi4800m;
wire cdxi5319m = cdxi4915m&r7m;
wire cdxi5320m = cdxi4743m&cdxi4920m;
wire cdxi5321m = cdxi4873m&r9m;
wire cdxi5322m = cdxi4916m&r13m;
wire cdxi5323m = cdxi4874m&r14m;
wire cdxi5324m = cdxi4875m&r18m;
wire cdxi5325m = cdxi4722m&r28m;
wire cdxi5326m = cdxi4711m&r29m;
wire cdxi5327m = cdxi4743m&r33m;
wire cdxi5328m = cdxi4712m&r43m;
wire cdxi5329m = (cdxi63m ^ cdxi5315m ^ cdxi5316m ^ cdxi5317m ^ cdxi5318m ^ cdxi5319m ^ cdxi5320m ^ cdxi5321m ^ cdxi5322m ^ cdxi5323m ^ cdxi5324m ^ cdxi5325m ^ cdxi5326m ^ cdxi5327m ^ cdxi5328m);
wire cdxi5330m = a1&cdxi5329m;
wire cdxi5331m = (reg_1_37);
wire cdxi5332m = (reg_1_71);
wire cdxi5333m = reg_1_2&cdxi4926m;
wire cdxi5334m = reg_1_1&cdxi5020m;
wire cdxi5335m = reg_1_1&cdxi5021m;
wire cdxi5336m = reg_1_1&cdxi5022m;
wire cdxi5337m = reg_1_3&reg_1_4&cdxi4884m;
wire cdxi5338m = reg_1_2&cdxi4929m;
wire cdxi5339m = reg_1_2&cdxi4930m;
wire cdxi5340m = reg_1_1&cdxi5023m;
wire cdxi5341m = reg_1_1&cdxi5024m;
wire cdxi5342m = reg_1_1&cdxi5025m;
wire cdxi5343m = reg_1_4&cdxi4886m;
wire cdxi5344m = reg_1_3&cdxi5331m;
wire cdxi5345m = reg_1_2&cdxi4925m;
wire cdxi5346m = reg_1_1&cdxi5019m;
wire cdxi5347m = (cdxi5333m ^ cdxi5334m ^ cdxi5335m ^ cdxi5336m ^ cdxi5337m ^ cdxi5338m ^ cdxi5339m ^ cdxi5340m ^ cdxi5341m ^ cdxi5342m ^ cdxi5343m ^ cdxi5344m ^ cdxi5345m ^ cdxi5346m ^ cdxi5332m);
wire cdxi5348m = reg_1_0&cdxi5347m;
wire cdxi5349m = cdxi4873m&cdxi4762m;
wire cdxi5350m = cdxi4874m&cdxi4762m;
wire cdxi5351m = cdxi4875m&cdxi4762m;
wire cdxi5352m = cdxi5349m&r0m;
wire cdxi5353m = cdxi5350m&r1m;
wire cdxi5354m = cdxi4875m&cdxi4826m;
wire cdxi5355m = cdxi4875m&cdxi4827m;
wire cdxi5356m = cdxi5083m&r7m;
wire cdxi5357m = cdxi5028m&r8m;
wire cdxi5358m = cdxi4873m&r10m;
wire cdxi5359m = cdxi4954m&r13m;
wire cdxi5360m = cdxi4874m&r15m;
wire cdxi5361m = cdxi4875m&r19m;
wire cdxi5362m = cdxi4762m&r28m;
wire cdxi5363m = cdxi4711m&r30m;
wire cdxi5364m = cdxi4743m&r34m;
wire cdxi5365m = cdxi4712m&r44m;
wire cdxi5366m = (cdxi64m ^ cdxi5352m ^ cdxi5353m ^ cdxi5354m ^ cdxi5355m ^ cdxi5356m ^ cdxi5357m ^ cdxi5358m ^ cdxi5359m ^ cdxi5360m ^ cdxi5361m ^ cdxi5362m ^ cdxi5363m ^ cdxi5364m ^ cdxi5365m);
wire cdxi5367m = a1&cdxi5366m;
wire cdxi5368m = (reg_1_38);
wire cdxi5369m = (reg_1_42);
wire cdxi5370m = (reg_1_72);
wire cdxi5371m = reg_1_2&reg_1_3&reg_1_5&cdxi4664m;
wire cdxi5372m = reg_1_1&cdxi5181m;
wire cdxi5373m = reg_1_1&cdxi5182m;
wire cdxi5374m = reg_1_1&cdxi5183m;
wire cdxi5375m = reg_1_3&reg_1_5&cdxi4884m;
wire cdxi5376m = reg_1_2&reg_1_5&cdxi4717m;
wire cdxi5377m = reg_1_2&reg_1_3&cdxi4963m;
wire cdxi5378m = reg_1_1&cdxi5184m;
wire cdxi5379m = reg_1_1&cdxi5185m;
wire cdxi5380m = reg_1_1&cdxi5186m;
wire cdxi5381m = reg_1_5&cdxi4886m;
wire cdxi5382m = reg_1_3&cdxi5368m;
wire cdxi5383m = reg_1_2&cdxi5369m;
wire cdxi5384m = reg_1_1&cdxi5180m;
wire cdxi5385m = (cdxi5371m ^ cdxi5372m ^ cdxi5373m ^ cdxi5374m ^ cdxi5375m ^ cdxi5376m ^ cdxi5377m ^ cdxi5378m ^ cdxi5379m ^ cdxi5380m ^ cdxi5381m ^ cdxi5382m ^ cdxi5383m ^ cdxi5384m ^ cdxi5370m);
wire cdxi5386m = reg_1_0&cdxi5385m;
wire cdxi5387m = cdxi4873m&cdxi4742m;
wire cdxi5388m = cdxi4874m&cdxi4742m;
wire cdxi5389m = cdxi4875m&cdxi4742m;
wire cdxi5390m = cdxi5387m&r0m;
wire cdxi5391m = cdxi4874m&cdxi4744m;
wire cdxi5392m = cdxi4875m&cdxi4808m;
wire cdxi5393m = cdxi4875m&cdxi4809m;
wire cdxi5394m = cdxi4711m&cdxi4900m;
wire cdxi5395m = cdxi4895m&r8m;
wire cdxi5396m = cdxi4873m&r11m;
wire cdxi5397m = cdxi4896m&r13m;
wire cdxi5398m = cdxi4874m&r16m;
wire cdxi5399m = cdxi4875m&r20m;
wire cdxi5400m = cdxi4742m&r28m;
wire cdxi5401m = cdxi4711m&r31m;
wire cdxi5402m = cdxi4743m&r35m;
wire cdxi5403m = cdxi4712m&r45m;
wire cdxi5404m = (cdxi65m ^ cdxi5390m ^ cdxi5391m ^ cdxi5392m ^ cdxi5393m ^ cdxi5394m ^ cdxi5395m ^ cdxi5396m ^ cdxi5397m ^ cdxi5398m ^ cdxi5399m ^ cdxi5400m ^ cdxi5401m ^ cdxi5402m ^ cdxi5403m);
wire cdxi5405m = a1&cdxi5404m;
wire cdxi5406m = (reg_1_43);
wire cdxi5407m = (reg_1_73);
wire cdxi5408m = reg_1_2&reg_1_3&reg_1_6&cdxi4664m;
wire cdxi5409m = reg_1_1&cdxi5198m;
wire cdxi5410m = reg_1_1&cdxi5199m;
wire cdxi5411m = reg_1_1&cdxi5200m;
wire cdxi5412m = reg_1_3&cdxi4910m;
wire cdxi5413m = reg_1_2&reg_1_6&cdxi4717m;
wire cdxi5414m = reg_1_2&reg_1_3&cdxi4905m;
wire cdxi5415m = reg_1_1&cdxi5201m;
wire cdxi5416m = reg_1_1&cdxi5202m;
wire cdxi5417m = reg_1_1&cdxi5203m;
wire cdxi5418m = reg_1_6&cdxi4886m;
wire cdxi5419m = reg_1_3&cdxi4906m;
wire cdxi5420m = reg_1_2&cdxi5406m;
wire cdxi5421m = reg_1_1&cdxi5197m;
wire cdxi5422m = (cdxi5408m ^ cdxi5409m ^ cdxi5410m ^ cdxi5411m ^ cdxi5412m ^ cdxi5413m ^ cdxi5414m ^ cdxi5415m ^ cdxi5416m ^ cdxi5417m ^ cdxi5418m ^ cdxi5419m ^ cdxi5420m ^ cdxi5421m ^ cdxi5407m);
wire cdxi5423m = reg_1_0&cdxi5422m;
wire cdxi5424m = cdxi4873m&cdxi4732m;
wire cdxi5425m = cdxi4874m&cdxi4732m;
wire cdxi5426m = cdxi4875m&cdxi4732m;
wire cdxi5427m = cdxi4873m&cdxi4733m;
wire cdxi5428m = cdxi4874m&cdxi4790m;
wire cdxi5429m = cdxi4875m&cdxi4753m;
wire cdxi5430m = cdxi4875m&cdxi4754m;
wire cdxi5431m = cdxi4934m&r7m;
wire cdxi5432m = cdxi4743m&cdxi4939m;
wire cdxi5433m = cdxi4873m&r12m;
wire cdxi5434m = cdxi4935m&r13m;
wire cdxi5435m = cdxi4874m&r17m;
wire cdxi5436m = cdxi4875m&r21m;
wire cdxi5437m = cdxi4732m&r28m;
wire cdxi5438m = cdxi4711m&r32m;
wire cdxi5439m = cdxi4743m&r36m;
wire cdxi5440m = cdxi4712m&r46m;
wire cdxi5441m = (cdxi66m ^ cdxi5427m ^ cdxi5428m ^ cdxi5429m ^ cdxi5430m ^ cdxi5431m ^ cdxi5432m ^ cdxi5433m ^ cdxi5434m ^ cdxi5435m ^ cdxi5436m ^ cdxi5437m ^ cdxi5438m ^ cdxi5439m ^ cdxi5440m);
wire cdxi5442m = a1&cdxi5441m;
wire cdxi5443m = (reg_1_40);
wire cdxi5444m = (reg_1_54);
wire cdxi5445m = (reg_1_74);
wire cdxi5446m = reg_1_2&cdxi4945m;
wire cdxi5447m = reg_1_1&reg_1_3&cdxi4795m;
wire cdxi5448m = reg_1_1&reg_1_2&cdxi4758m;
wire cdxi5449m = reg_1_1&reg_1_2&cdxi4759m;
wire cdxi5450m = reg_1_3&reg_1_7&cdxi4884m;
wire cdxi5451m = reg_1_2&cdxi4948m;
wire cdxi5452m = reg_1_2&cdxi4949m;
wire cdxi5453m = reg_1_1&reg_1_7&cdxi4885m;
wire cdxi5454m = reg_1_1&reg_1_3&cdxi4794m;
wire cdxi5455m = reg_1_1&reg_1_2&cdxi4757m;
wire cdxi5456m = reg_1_7&cdxi4886m;
wire cdxi5457m = reg_1_3&cdxi5443m;
wire cdxi5458m = reg_1_2&cdxi4944m;
wire cdxi5459m = reg_1_1&cdxi5444m;
wire cdxi5460m = (cdxi5446m ^ cdxi5447m ^ cdxi5448m ^ cdxi5449m ^ cdxi5450m ^ cdxi5451m ^ cdxi5452m ^ cdxi5453m ^ cdxi5454m ^ cdxi5455m ^ cdxi5456m ^ cdxi5457m ^ cdxi5458m ^ cdxi5459m ^ cdxi5445m);
wire cdxi5461m = reg_1_0&cdxi5460m;
wire cdxi5462m = cdxi4743m&cdxi4973m;
wire cdxi5463m = cdxi4916m&cdxi4742m;
wire cdxi5464m = cdxi4743m&cdxi4974m;
wire cdxi5465m = cdxi4916m&cdxi4744m;
wire cdxi5466m = cdxi4875m&cdxi4817m;
wire cdxi5467m = cdxi4875m&cdxi4818m;
wire cdxi5468m = cdxi4722m&cdxi4900m;
wire cdxi5469m = cdxi4895m&r9m;
wire cdxi5470m = cdxi4743m&cdxi4978m;
wire cdxi5471m = cdxi4896m&r14m;
wire cdxi5472m = cdxi4916m&r16m;
wire cdxi5473m = cdxi4875m&r23m;
wire cdxi5474m = cdxi4742m&r29m;
wire cdxi5475m = cdxi4722m&r31m;
wire cdxi5476m = cdxi4743m&r38m;
wire cdxi5477m = cdxi4712m&r48m;
wire cdxi5478m = (cdxi68m ^ cdxi5464m ^ cdxi5465m ^ cdxi5466m ^ cdxi5467m ^ cdxi5468m ^ cdxi5469m ^ cdxi5470m ^ cdxi5471m ^ cdxi5472m ^ cdxi5473m ^ cdxi5474m ^ cdxi5475m ^ cdxi5476m ^ cdxi5477m);
wire cdxi5479m = a1&cdxi5478m;
wire cdxi5480m = (reg_1_76);
wire cdxi5481m = reg_1_2&cdxi4983m;
wire cdxi5482m = reg_1_1&cdxi5056m;
wire cdxi5483m = reg_1_1&cdxi5057m;
wire cdxi5484m = reg_1_1&cdxi5058m;
wire cdxi5485m = reg_1_4&cdxi4910m;
wire cdxi5486m = reg_1_2&cdxi4986m;
wire cdxi5487m = reg_1_2&cdxi4987m;
wire cdxi5488m = reg_1_1&cdxi5059m;
wire cdxi5489m = reg_1_1&cdxi5060m;
wire cdxi5490m = reg_1_1&cdxi5061m;
wire cdxi5491m = reg_1_6&cdxi5331m;
wire cdxi5492m = reg_1_4&cdxi4906m;
wire cdxi5493m = reg_1_2&cdxi4982m;
wire cdxi5494m = reg_1_1&cdxi5055m;
wire cdxi5495m = (cdxi5481m ^ cdxi5482m ^ cdxi5483m ^ cdxi5484m ^ cdxi5485m ^ cdxi5486m ^ cdxi5487m ^ cdxi5488m ^ cdxi5489m ^ cdxi5490m ^ cdxi5491m ^ cdxi5492m ^ cdxi5493m ^ cdxi5494m ^ cdxi5480m);
wire cdxi5496m = reg_1_0&cdxi5495m;
wire cdxi5497m = cdxi5028m&cdxi4742m;
wire cdxi5498m = cdxi4954m&cdxi4742m;
wire cdxi5499m = cdxi5497m&r0m;
wire cdxi5500m = cdxi4954m&cdxi4744m;
wire cdxi5501m = cdxi4875m&cdxi4772m;
wire cdxi5502m = cdxi4875m&cdxi4773m;
wire cdxi5503m = cdxi4762m&cdxi4900m;
wire cdxi5504m = cdxi4895m&r10m;
wire cdxi5505m = cdxi5028m&r11m;
wire cdxi5506m = cdxi4896m&r15m;
wire cdxi5507m = cdxi4954m&r16m;
wire cdxi5508m = cdxi4875m&r25m;
wire cdxi5509m = cdxi4742m&r30m;
wire cdxi5510m = cdxi4762m&r31m;
wire cdxi5511m = cdxi4743m&r40m;
wire cdxi5512m = cdxi4712m&r50m;
wire cdxi5513m = (cdxi70m ^ cdxi5499m ^ cdxi5500m ^ cdxi5501m ^ cdxi5502m ^ cdxi5503m ^ cdxi5504m ^ cdxi5505m ^ cdxi5506m ^ cdxi5507m ^ cdxi5508m ^ cdxi5509m ^ cdxi5510m ^ cdxi5511m ^ cdxi5512m);
wire cdxi5514m = a1&cdxi5513m;
wire cdxi5515m = (reg_1_48);
wire cdxi5516m = (reg_1_78);
wire cdxi5517m = reg_1_2&reg_1_5&reg_1_6&cdxi4664m;
wire cdxi5518m = reg_1_1&cdxi5219m;
wire cdxi5519m = reg_1_1&cdxi5220m;
wire cdxi5520m = reg_1_1&cdxi5221m;
wire cdxi5521m = reg_1_5&cdxi4910m;
wire cdxi5522m = reg_1_2&reg_1_6&cdxi4963m;
wire cdxi5523m = reg_1_2&reg_1_5&cdxi4905m;
wire cdxi5524m = reg_1_1&cdxi5222m;
wire cdxi5525m = reg_1_1&cdxi5223m;
wire cdxi5526m = reg_1_1&cdxi5224m;
wire cdxi5527m = reg_1_6&cdxi5368m;
wire cdxi5528m = reg_1_5&cdxi4906m;
wire cdxi5529m = reg_1_2&cdxi5515m;
wire cdxi5530m = reg_1_1&cdxi5218m;
wire cdxi5531m = (cdxi5517m ^ cdxi5518m ^ cdxi5519m ^ cdxi5520m ^ cdxi5521m ^ cdxi5522m ^ cdxi5523m ^ cdxi5524m ^ cdxi5525m ^ cdxi5526m ^ cdxi5527m ^ cdxi5528m ^ cdxi5529m ^ cdxi5530m ^ cdxi5516m);
wire cdxi5532m = reg_1_0&cdxi5531m;
wire cdxi5533m = cdxi4895m&cdxi4732m;
wire cdxi5534m = cdxi4896m&cdxi4732m;
wire cdxi5535m = cdxi4895m&cdxi4733m;
wire cdxi5536m = cdxi4896m&cdxi4790m;
wire cdxi5537m = cdxi4875m&cdxi4850m;
wire cdxi5538m = cdxi4875m&cdxi4851m;
wire cdxi5539m = cdxi5154m&r7m;
wire cdxi5540m = cdxi5065m&r11m;
wire cdxi5541m = cdxi4895m&r12m;
wire cdxi5542m = cdxi4935m&r16m;
wire cdxi5543m = cdxi4896m&r17m;
wire cdxi5544m = cdxi4875m&r27m;
wire cdxi5545m = cdxi4732m&r31m;
wire cdxi5546m = cdxi4742m&r32m;
wire cdxi5547m = cdxi4743m&r42m;
wire cdxi5548m = cdxi4712m&r52m;
wire cdxi5549m = (cdxi72m ^ cdxi5535m ^ cdxi5536m ^ cdxi5537m ^ cdxi5538m ^ cdxi5539m ^ cdxi5540m ^ cdxi5541m ^ cdxi5542m ^ cdxi5543m ^ cdxi5544m ^ cdxi5545m ^ cdxi5546m ^ cdxi5547m ^ cdxi5548m);
wire cdxi5550m = a1&cdxi5549m;
wire cdxi5551m = (reg_1_50);
wire cdxi5552m = (reg_1_60);
wire cdxi5553m = (reg_1_80);
wire cdxi5554m = reg_1_2&reg_1_6&cdxi4738m;
wire cdxi5555m = reg_1_1&reg_1_6&cdxi4795m;
wire cdxi5556m = reg_1_1&reg_1_2&cdxi4855m;
wire cdxi5557m = reg_1_1&reg_1_2&cdxi4856m;
wire cdxi5558m = reg_1_6&reg_1_7&cdxi4884m;
wire cdxi5559m = reg_1_2&reg_1_7&cdxi4905m;
wire cdxi5560m = reg_1_2&reg_1_6&cdxi4737m;
wire cdxi5561m = reg_1_1&reg_1_7&cdxi4748m;
wire cdxi5562m = reg_1_1&reg_1_6&cdxi4794m;
wire cdxi5563m = reg_1_1&reg_1_2&cdxi4854m;
wire cdxi5564m = reg_1_7&cdxi4906m;
wire cdxi5565m = reg_1_6&cdxi5443m;
wire cdxi5566m = reg_1_2&cdxi5551m;
wire cdxi5567m = reg_1_1&cdxi5552m;
wire cdxi5568m = (cdxi5554m ^ cdxi5555m ^ cdxi5556m ^ cdxi5557m ^ cdxi5558m ^ cdxi5559m ^ cdxi5560m ^ cdxi5561m ^ cdxi5562m ^ cdxi5563m ^ cdxi5564m ^ cdxi5565m ^ cdxi5566m ^ cdxi5567m ^ cdxi5553m);
wire cdxi5569m = reg_1_0&cdxi5568m;
wire cdxi5570m = cdxi4915m&cdxi4742m;
wire cdxi5571m = cdxi5570m&r0m;
wire cdxi5572m = cdxi4916m&cdxi4808m;
wire cdxi5573m = cdxi4874m&cdxi4817m;
wire cdxi5574m = cdxi4874m&cdxi4818m;
wire cdxi5575m = cdxi4973m&r8m;
wire cdxi5576m = cdxi4711m&cdxi4977m;
wire cdxi5577m = cdxi4915m&r11m;
wire cdxi5578m = cdxi4896m&r18m;
wire cdxi5579m = cdxi4916m&r20m;
wire cdxi5580m = cdxi4874m&r23m;
wire cdxi5581m = cdxi4742m&r33m;
wire cdxi5582m = cdxi4722m&r35m;
wire cdxi5583m = cdxi4711m&r38m;
wire cdxi5584m = cdxi4712m&r54m;
wire cdxi5585m = (cdxi74m ^ cdxi5571m ^ cdxi5572m ^ cdxi5573m ^ cdxi5574m ^ cdxi5575m ^ cdxi5576m ^ cdxi5577m ^ cdxi5578m ^ cdxi5579m ^ cdxi5580m ^ cdxi5581m ^ cdxi5582m ^ cdxi5583m ^ cdxi5584m);
wire cdxi5586m = a1&cdxi5585m;
wire cdxi5587m = (reg_1_82);
wire cdxi5588m = reg_1_3&cdxi4983m;
wire cdxi5589m = reg_1_1&cdxi5111m;
wire cdxi5590m = reg_1_1&cdxi5112m;
wire cdxi5591m = reg_1_1&cdxi5113m;
wire cdxi5592m = reg_1_4&reg_1_6&cdxi4717m;
wire cdxi5593m = reg_1_3&cdxi4986m;
wire cdxi5594m = reg_1_3&cdxi4987m;
wire cdxi5595m = reg_1_1&cdxi5114m;
wire cdxi5596m = reg_1_1&cdxi5115m;
wire cdxi5597m = reg_1_1&cdxi5116m;
wire cdxi5598m = reg_1_6&cdxi4925m;
wire cdxi5599m = reg_1_4&cdxi5406m;
wire cdxi5600m = reg_1_3&cdxi4982m;
wire cdxi5601m = reg_1_1&cdxi5110m;
wire cdxi5602m = (cdxi5588m ^ cdxi5589m ^ cdxi5590m ^ cdxi5591m ^ cdxi5592m ^ cdxi5593m ^ cdxi5594m ^ cdxi5595m ^ cdxi5596m ^ cdxi5597m ^ cdxi5598m ^ cdxi5599m ^ cdxi5600m ^ cdxi5601m ^ cdxi5587m);
wire cdxi5603m = reg_1_0&cdxi5602m;
wire cdxi5604m = cdxi4915m&cdxi4732m;
wire cdxi5605m = cdxi4916m&cdxi4732m;
wire cdxi5606m = cdxi4915m&cdxi4733m;
wire cdxi5607m = cdxi4916m&cdxi4753m;
wire cdxi5608m = cdxi4874m&cdxi4839m;
wire cdxi5609m = cdxi4874m&cdxi4840m;
wire cdxi5610m = cdxi4722m&cdxi4939m;
wire cdxi5611m = cdxi4934m&r9m;
wire cdxi5612m = cdxi4915m&r12m;
wire cdxi5613m = cdxi4935m&r18m;
wire cdxi5614m = cdxi4916m&r21m;
wire cdxi5615m = cdxi4874m&r24m;
wire cdxi5616m = cdxi4732m&r33m;
wire cdxi5617m = cdxi4722m&r36m;
wire cdxi5618m = cdxi4711m&r39m;
wire cdxi5619m = cdxi4712m&r55m;
wire cdxi5620m = (cdxi75m ^ cdxi5606m ^ cdxi5607m ^ cdxi5608m ^ cdxi5609m ^ cdxi5610m ^ cdxi5611m ^ cdxi5612m ^ cdxi5613m ^ cdxi5614m ^ cdxi5615m ^ cdxi5616m ^ cdxi5617m ^ cdxi5618m ^ cdxi5619m);
wire cdxi5621m = a1&cdxi5620m;
wire cdxi5622m = (reg_1_47);
wire cdxi5623m = (reg_1_83);
wire cdxi5624m = reg_1_3&reg_1_4&cdxi4738m;
wire cdxi5625m = reg_1_1&cdxi5278m;
wire cdxi5626m = reg_1_1&cdxi5279m;
wire cdxi5627m = reg_1_1&cdxi5280m;
wire cdxi5628m = reg_1_4&cdxi4948m;
wire cdxi5629m = reg_1_3&reg_1_7&cdxi4727m;
wire cdxi5630m = reg_1_3&reg_1_4&cdxi4737m;
wire cdxi5631m = reg_1_1&cdxi5281m;
wire cdxi5632m = reg_1_1&cdxi5282m;
wire cdxi5633m = reg_1_1&cdxi5283m;
wire cdxi5634m = reg_1_7&cdxi4925m;
wire cdxi5635m = reg_1_4&cdxi4944m;
wire cdxi5636m = reg_1_3&cdxi5622m;
wire cdxi5637m = reg_1_1&cdxi5277m;
wire cdxi5638m = (cdxi5624m ^ cdxi5625m ^ cdxi5626m ^ cdxi5627m ^ cdxi5628m ^ cdxi5629m ^ cdxi5630m ^ cdxi5631m ^ cdxi5632m ^ cdxi5633m ^ cdxi5634m ^ cdxi5635m ^ cdxi5636m ^ cdxi5637m ^ cdxi5623m);
wire cdxi5639m = reg_1_0&cdxi5638m;
wire cdxi5640m = cdxi4711m&cdxi4991m;
wire cdxi5641m = cdxi4954m&cdxi4732m;
wire cdxi5642m = cdxi4711m&cdxi4992m;
wire cdxi5643m = cdxi4954m&cdxi4753m;
wire cdxi5644m = cdxi4874m&cdxi4781m;
wire cdxi5645m = cdxi4874m&cdxi4782m;
wire cdxi5646m = cdxi4762m&cdxi4939m;
wire cdxi5647m = cdxi4934m&r10m;
wire cdxi5648m = cdxi4711m&cdxi4996m;
wire cdxi5649m = cdxi4935m&r19m;
wire cdxi5650m = cdxi4954m&r21m;
wire cdxi5651m = cdxi4874m&r26m;
wire cdxi5652m = cdxi4732m&r34m;
wire cdxi5653m = cdxi4762m&r36m;
wire cdxi5654m = cdxi4711m&r41m;
wire cdxi5655m = cdxi4712m&r57m;
wire cdxi5656m = (cdxi77m ^ cdxi5642m ^ cdxi5643m ^ cdxi5644m ^ cdxi5645m ^ cdxi5646m ^ cdxi5647m ^ cdxi5648m ^ cdxi5649m ^ cdxi5650m ^ cdxi5651m ^ cdxi5652m ^ cdxi5653m ^ cdxi5654m ^ cdxi5655m);
wire cdxi5657m = a1&cdxi5656m;
wire cdxi5658m = (reg_1_85);
wire cdxi5659m = reg_1_3&cdxi5001m;
wire cdxi5660m = reg_1_1&cdxi5128m;
wire cdxi5661m = reg_1_1&cdxi5129m;
wire cdxi5662m = reg_1_1&cdxi5130m;
wire cdxi5663m = reg_1_5&cdxi4948m;
wire cdxi5664m = reg_1_3&cdxi5004m;
wire cdxi5665m = reg_1_3&cdxi5005m;
wire cdxi5666m = reg_1_1&cdxi5131m;
wire cdxi5667m = reg_1_1&cdxi5132m;
wire cdxi5668m = reg_1_1&cdxi5133m;
wire cdxi5669m = reg_1_7&cdxi5369m;
wire cdxi5670m = reg_1_5&cdxi4944m;
wire cdxi5671m = reg_1_3&cdxi5000m;
wire cdxi5672m = reg_1_1&cdxi5127m;
wire cdxi5673m = (cdxi5659m ^ cdxi5660m ^ cdxi5661m ^ cdxi5662m ^ cdxi5663m ^ cdxi5664m ^ cdxi5665m ^ cdxi5666m ^ cdxi5667m ^ cdxi5668m ^ cdxi5669m ^ cdxi5670m ^ cdxi5671m ^ cdxi5672m ^ cdxi5658m);
wire cdxi5674m = reg_1_0&cdxi5673m;
wire cdxi5675m = cdxi5101m&cdxi4732m;
wire cdxi5676m = cdxi5101m&cdxi4733m;
wire cdxi5677m = cdxi4896m&cdxi4753m;
wire cdxi5678m = cdxi4874m&cdxi4850m;
wire cdxi5679m = cdxi4874m&cdxi4851m;
wire cdxi5680m = cdxi4742m&cdxi4939m;
wire cdxi5681m = cdxi4934m&r11m;
wire cdxi5682m = cdxi5101m&r12m;
wire cdxi5683m = cdxi4935m&r20m;
wire cdxi5684m = cdxi4896m&r21m;
wire cdxi5685m = cdxi4874m&r27m;
wire cdxi5686m = cdxi4732m&r35m;
wire cdxi5687m = cdxi4742m&r36m;
wire cdxi5688m = cdxi4711m&r42m;
wire cdxi5689m = cdxi4712m&r58m;
wire cdxi5690m = (cdxi78m ^ cdxi5676m ^ cdxi5677m ^ cdxi5678m ^ cdxi5679m ^ cdxi5680m ^ cdxi5681m ^ cdxi5682m ^ cdxi5683m ^ cdxi5684m ^ cdxi5685m ^ cdxi5686m ^ cdxi5687m ^ cdxi5688m ^ cdxi5689m);
wire cdxi5691m = a1&cdxi5690m;
wire cdxi5692m = (reg_1_66);
wire cdxi5693m = (reg_1_86);
wire cdxi5694m = reg_1_3&reg_1_6&cdxi4738m;
wire cdxi5695m = reg_1_1&reg_1_6&cdxi4758m;
wire cdxi5696m = reg_1_1&reg_1_3&cdxi4855m;
wire cdxi5697m = reg_1_1&reg_1_3&cdxi4856m;
wire cdxi5698m = reg_1_6&cdxi4948m;
wire cdxi5699m = reg_1_3&reg_1_7&cdxi4905m;
wire cdxi5700m = reg_1_3&reg_1_6&cdxi4737m;
wire cdxi5701m = reg_1_1&reg_1_7&cdxi4812m;
wire cdxi5702m = reg_1_1&reg_1_6&cdxi4757m;
wire cdxi5703m = reg_1_1&reg_1_3&cdxi4854m;
wire cdxi5704m = reg_1_7&cdxi5406m;
wire cdxi5705m = reg_1_6&cdxi4944m;
wire cdxi5706m = reg_1_3&cdxi5551m;
wire cdxi5707m = reg_1_1&cdxi5692m;
wire cdxi5708m = (cdxi5694m ^ cdxi5695m ^ cdxi5696m ^ cdxi5697m ^ cdxi5698m ^ cdxi5699m ^ cdxi5700m ^ cdxi5701m ^ cdxi5702m ^ cdxi5703m ^ cdxi5704m ^ cdxi5705m ^ cdxi5706m ^ cdxi5707m ^ cdxi5693m);
wire cdxi5709m = reg_1_0&cdxi5708m;
wire cdxi5710m = cdxi4953m&cdxi4732m;
wire cdxi5711m = cdxi4916m&cdxi4762m;
wire cdxi5712m = cdxi4953m&cdxi4733m;
wire cdxi5713m = cdxi4954m&cdxi4839m;
wire cdxi5714m = cdxi4916m&cdxi4781m;
wire cdxi5715m = cdxi4916m&cdxi4782m;
wire cdxi5716m = cdxi4991m&r9m;
wire cdxi5717m = cdxi4722m&cdxi4995m;
wire cdxi5718m = cdxi4953m&r12m;
wire cdxi5719m = cdxi4935m&r22m;
wire cdxi5720m = cdxi4954m&r24m;
wire cdxi5721m = cdxi4916m&r26m;
wire cdxi5722m = cdxi4732m&r37m;
wire cdxi5723m = cdxi4762m&r39m;
wire cdxi5724m = cdxi4722m&r41m;
wire cdxi5725m = cdxi4712m&r60m;
wire cdxi5726m = (cdxi80m ^ cdxi5712m ^ cdxi5713m ^ cdxi5714m ^ cdxi5715m ^ cdxi5716m ^ cdxi5717m ^ cdxi5718m ^ cdxi5719m ^ cdxi5720m ^ cdxi5721m ^ cdxi5722m ^ cdxi5723m ^ cdxi5724m ^ cdxi5725m);
wire cdxi5727m = a1&cdxi5726m;
wire cdxi5728m = (reg_1_88);
wire cdxi5729m = reg_1_4&cdxi5001m;
wire cdxi5730m = reg_1_1&cdxi5301m;
wire cdxi5731m = reg_1_1&cdxi5302m;
wire cdxi5732m = reg_1_1&cdxi5303m;
wire cdxi5733m = reg_1_5&reg_1_7&cdxi4727m;
wire cdxi5734m = reg_1_4&cdxi5004m;
wire cdxi5735m = reg_1_4&cdxi5005m;
wire cdxi5736m = reg_1_1&cdxi5304m;
wire cdxi5737m = reg_1_1&cdxi5305m;
wire cdxi5738m = reg_1_1&cdxi5306m;
wire cdxi5739m = reg_1_7&cdxi4964m;
wire cdxi5740m = reg_1_5&cdxi5622m;
wire cdxi5741m = reg_1_4&cdxi5000m;
wire cdxi5742m = reg_1_1&cdxi5300m;
wire cdxi5743m = (cdxi5729m ^ cdxi5730m ^ cdxi5731m ^ cdxi5732m ^ cdxi5733m ^ cdxi5734m ^ cdxi5735m ^ cdxi5736m ^ cdxi5737m ^ cdxi5738m ^ cdxi5739m ^ cdxi5740m ^ cdxi5741m ^ cdxi5742m ^ cdxi5728m);
wire cdxi5744m = reg_1_0&cdxi5743m;
wire cdxi5745m = cdxi4973m&cdxi4732m;
wire cdxi5746m = cdxi4973m&cdxi4733m;
wire cdxi5747m = cdxi4896m&cdxi4839m;
wire cdxi5748m = cdxi4916m&cdxi4850m;
wire cdxi5749m = cdxi4916m&cdxi4851m;
wire cdxi5750m = cdxi5154m&r9m;
wire cdxi5751m = cdxi5064m&r11m;
wire cdxi5752m = cdxi4973m&r12m;
wire cdxi5753m = cdxi4935m&r23m;
wire cdxi5754m = cdxi4896m&r24m;
wire cdxi5755m = cdxi4916m&r27m;
wire cdxi5756m = cdxi4732m&r38m;
wire cdxi5757m = cdxi4742m&r39m;
wire cdxi5758m = cdxi4722m&r42m;
wire cdxi5759m = cdxi4712m&r61m;
wire cdxi5760m = (cdxi81m ^ cdxi5746m ^ cdxi5747m ^ cdxi5748m ^ cdxi5749m ^ cdxi5750m ^ cdxi5751m ^ cdxi5752m ^ cdxi5753m ^ cdxi5754m ^ cdxi5755m ^ cdxi5756m ^ cdxi5757m ^ cdxi5758m ^ cdxi5759m);
wire cdxi5761m = a1&cdxi5760m;
wire cdxi5762m = (reg_1_89);
wire cdxi5763m = reg_1_4&reg_1_6&cdxi4738m;
wire cdxi5764m = reg_1_1&cdxi5259m;
wire cdxi5765m = reg_1_1&cdxi5260m;
wire cdxi5766m = reg_1_1&cdxi5261m;
wire cdxi5767m = reg_1_6&reg_1_7&cdxi4727m;
wire cdxi5768m = reg_1_4&reg_1_7&cdxi4905m;
wire cdxi5769m = reg_1_4&reg_1_6&cdxi4737m;
wire cdxi5770m = reg_1_1&cdxi5262m;
wire cdxi5771m = reg_1_1&cdxi5263m;
wire cdxi5772m = reg_1_1&cdxi5264m;
wire cdxi5773m = reg_1_7&cdxi4982m;
wire cdxi5774m = reg_1_6&cdxi5622m;
wire cdxi5775m = reg_1_4&cdxi5551m;
wire cdxi5776m = reg_1_1&cdxi5258m;
wire cdxi5777m = (cdxi5763m ^ cdxi5764m ^ cdxi5765m ^ cdxi5766m ^ cdxi5767m ^ cdxi5768m ^ cdxi5769m ^ cdxi5770m ^ cdxi5771m ^ cdxi5772m ^ cdxi5773m ^ cdxi5774m ^ cdxi5775m ^ cdxi5776m ^ cdxi5762m);
wire cdxi5778m = reg_1_0&cdxi5777m;
wire cdxi5779m = cdxi4915m&cdxi4762m;
wire cdxi5780m = cdxi4743m&cdxi4953m;
wire cdxi5781m = cdxi5779m&r1m;
wire cdxi5782m = cdxi5009m&cdxi4826m;
wire cdxi5783m = cdxi4873m&cdxi4763m;
wire cdxi5784m = cdxi4873m&cdxi4764m;
wire cdxi5785m = cdxi4953m&r13m;
wire cdxi5786m = cdxi4711m&cdxi5032m;
wire cdxi5787m = cdxi4915m&r15m;
wire cdxi5788m = cdxi5028m&r18m;
wire cdxi5789m = cdxi5009m&r19m;
wire cdxi5790m = cdxi4873m&r22m;
wire cdxi5791m = cdxi4762m&r43m;
wire cdxi5792m = cdxi4722m&r44m;
wire cdxi5793m = cdxi4711m&r47m;
wire cdxi5794m = cdxi4743m&r53m;
wire cdxi5795m = (cdxi83m ^ cdxi5781m ^ cdxi5782m ^ cdxi5783m ^ cdxi5784m ^ cdxi5785m ^ cdxi5786m ^ cdxi5787m ^ cdxi5788m ^ cdxi5789m ^ cdxi5790m ^ cdxi5791m ^ cdxi5792m ^ cdxi5793m ^ cdxi5794m);
wire cdxi5796m = a1&cdxi5795m;
wire cdxi5797m = (reg_1_91);
wire cdxi5798m = reg_1_3&cdxi5039m;
wire cdxi5799m = reg_1_2&cdxi5093m;
wire cdxi5800m = reg_1_2&cdxi5094m;
wire cdxi5801m = reg_1_2&cdxi5095m;
wire cdxi5802m = reg_1_4&cdxi5184m;
wire cdxi5803m = reg_1_3&cdxi5042m;
wire cdxi5804m = reg_1_3&cdxi5043m;
wire cdxi5805m = reg_1_2&cdxi5096m;
wire cdxi5806m = reg_1_2&cdxi5097m;
wire cdxi5807m = reg_1_2&cdxi5098m;
wire cdxi5808m = reg_1_5&cdxi5019m;
wire cdxi5809m = reg_1_4&cdxi5180m;
wire cdxi5810m = reg_1_3&cdxi5038m;
wire cdxi5811m = reg_1_2&cdxi5092m;
wire cdxi5812m = (cdxi5798m ^ cdxi5799m ^ cdxi5800m ^ cdxi5801m ^ cdxi5802m ^ cdxi5803m ^ cdxi5804m ^ cdxi5805m ^ cdxi5806m ^ cdxi5807m ^ cdxi5808m ^ cdxi5809m ^ cdxi5810m ^ cdxi5811m ^ cdxi5797m);
wire cdxi5813m = reg_1_0&cdxi5812m;
wire cdxi5814m = cdxi5009m&cdxi4732m;
wire cdxi5815m = cdxi4915m&cdxi4790m;
wire cdxi5816m = cdxi5009m&cdxi4753m;
wire cdxi5817m = cdxi4873m&cdxi4839m;
wire cdxi5818m = cdxi4873m&cdxi4840m;
wire cdxi5819m = cdxi5064m&r13m;
wire cdxi5820m = cdxi4934m&r14m;
wire cdxi5821m = cdxi4915m&r17m;
wire cdxi5822m = cdxi5065m&r18m;
wire cdxi5823m = cdxi5009m&r21m;
wire cdxi5824m = cdxi4873m&r24m;
wire cdxi5825m = cdxi4732m&r43m;
wire cdxi5826m = cdxi4722m&r46m;
wire cdxi5827m = cdxi4711m&r49m;
wire cdxi5828m = cdxi4743m&r55m;
wire cdxi5829m = (cdxi85m ^ cdxi5815m ^ cdxi5816m ^ cdxi5817m ^ cdxi5818m ^ cdxi5819m ^ cdxi5820m ^ cdxi5821m ^ cdxi5822m ^ cdxi5823m ^ cdxi5824m ^ cdxi5825m ^ cdxi5826m ^ cdxi5827m ^ cdxi5828m);
wire cdxi5830m = a1&cdxi5829m;
wire cdxi5831m = (reg_1_93);
wire cdxi5832m = reg_1_3&cdxi5075m;
wire cdxi5833m = reg_1_2&cdxi5278m;
wire cdxi5834m = reg_1_2&cdxi5279m;
wire cdxi5835m = reg_1_2&cdxi5280m;
wire cdxi5836m = reg_1_4&reg_1_7&cdxi4885m;
wire cdxi5837m = reg_1_3&cdxi5078m;
wire cdxi5838m = reg_1_3&cdxi5079m;
wire cdxi5839m = reg_1_2&cdxi5281m;
wire cdxi5840m = reg_1_2&cdxi5282m;
wire cdxi5841m = reg_1_2&cdxi5283m;
wire cdxi5842m = reg_1_7&cdxi5019m;
wire cdxi5843m = reg_1_4&cdxi5444m;
wire cdxi5844m = reg_1_3&cdxi5074m;
wire cdxi5845m = reg_1_2&cdxi5277m;
wire cdxi5846m = (cdxi5832m ^ cdxi5833m ^ cdxi5834m ^ cdxi5835m ^ cdxi5836m ^ cdxi5837m ^ cdxi5838m ^ cdxi5839m ^ cdxi5840m ^ cdxi5841m ^ cdxi5842m ^ cdxi5843m ^ cdxi5844m ^ cdxi5845m ^ cdxi5831m);
wire cdxi5847m = reg_1_0&cdxi5846m;
wire cdxi5848m = cdxi5083m&cdxi4742m;
wire cdxi5849m = cdxi5083m&cdxi4744m;
wire cdxi5850m = cdxi5028m&cdxi4808m;
wire cdxi5851m = cdxi4873m&cdxi4772m;
wire cdxi5852m = cdxi4873m&cdxi4773m;
wire cdxi5853m = cdxi5136m&r13m;
wire cdxi5854m = cdxi5101m&r15m;
wire cdxi5855m = cdxi5083m&r16m;
wire cdxi5856m = cdxi4895m&r19m;
wire cdxi5857m = cdxi5028m&r20m;
wire cdxi5858m = cdxi4873m&r25m;
wire cdxi5859m = cdxi4742m&r44m;
wire cdxi5860m = cdxi4762m&r45m;
wire cdxi5861m = cdxi4711m&r50m;
wire cdxi5862m = cdxi4743m&r56m;
wire cdxi5863m = (cdxi86m ^ cdxi5849m ^ cdxi5850m ^ cdxi5851m ^ cdxi5852m ^ cdxi5853m ^ cdxi5854m ^ cdxi5855m ^ cdxi5856m ^ cdxi5857m ^ cdxi5858m ^ cdxi5859m ^ cdxi5860m ^ cdxi5861m ^ cdxi5862m);
wire cdxi5864m = a1&cdxi5863m;
wire cdxi5865m = (reg_1_64);
wire cdxi5866m = (reg_1_94);
wire cdxi5867m = reg_1_3&cdxi5219m;
wire cdxi5868m = reg_1_2&reg_1_5&cdxi4813m;
wire cdxi5869m = reg_1_2&reg_1_3&cdxi4777m;
wire cdxi5870m = reg_1_2&reg_1_3&cdxi4778m;
wire cdxi5871m = reg_1_5&cdxi5201m;
wire cdxi5872m = reg_1_3&cdxi5222m;
wire cdxi5873m = reg_1_3&cdxi5223m;
wire cdxi5874m = reg_1_2&reg_1_6&cdxi4830m;
wire cdxi5875m = reg_1_2&reg_1_5&cdxi4812m;
wire cdxi5876m = reg_1_2&reg_1_3&cdxi4776m;
wire cdxi5877m = reg_1_6&cdxi5180m;
wire cdxi5878m = reg_1_5&cdxi5197m;
wire cdxi5879m = reg_1_3&cdxi5218m;
wire cdxi5880m = reg_1_2&cdxi5865m;
wire cdxi5881m = (cdxi5867m ^ cdxi5868m ^ cdxi5869m ^ cdxi5870m ^ cdxi5871m ^ cdxi5872m ^ cdxi5873m ^ cdxi5874m ^ cdxi5875m ^ cdxi5876m ^ cdxi5877m ^ cdxi5878m ^ cdxi5879m ^ cdxi5880m ^ cdxi5866m);
wire cdxi5882m = reg_1_0&cdxi5881m;
wire cdxi5883m = cdxi4743m&cdxi4991m;
wire cdxi5884m = cdxi5083m&cdxi4790m;
wire cdxi5885m = cdxi5028m&cdxi4753m;
wire cdxi5886m = cdxi4873m&cdxi4781m;
wire cdxi5887m = cdxi4873m&cdxi4782m;
wire cdxi5888m = cdxi4991m&r13m;
wire cdxi5889m = cdxi4934m&r15m;
wire cdxi5890m = cdxi5083m&r17m;
wire cdxi5891m = cdxi5065m&r19m;
wire cdxi5892m = cdxi5028m&r21m;
wire cdxi5893m = cdxi4873m&r26m;
wire cdxi5894m = cdxi4732m&r44m;
wire cdxi5895m = cdxi4762m&r46m;
wire cdxi5896m = cdxi4711m&r51m;
wire cdxi5897m = cdxi4743m&r57m;
wire cdxi5898m = (cdxi87m ^ cdxi5884m ^ cdxi5885m ^ cdxi5886m ^ cdxi5887m ^ cdxi5888m ^ cdxi5889m ^ cdxi5890m ^ cdxi5891m ^ cdxi5892m ^ cdxi5893m ^ cdxi5894m ^ cdxi5895m ^ cdxi5896m ^ cdxi5897m);
wire cdxi5899m = a1&cdxi5898m;
wire cdxi5900m = (reg_1_95);
wire cdxi5901m = reg_1_3&cdxi5236m;
wire cdxi5902m = reg_1_2&cdxi5128m;
wire cdxi5903m = reg_1_2&cdxi5129m;
wire cdxi5904m = reg_1_2&cdxi5130m;
wire cdxi5905m = reg_1_5&reg_1_7&cdxi4885m;
wire cdxi5906m = reg_1_3&cdxi5239m;
wire cdxi5907m = reg_1_3&cdxi5240m;
wire cdxi5908m = reg_1_2&cdxi5131m;
wire cdxi5909m = reg_1_2&cdxi5132m;
wire cdxi5910m = reg_1_2&cdxi5133m;
wire cdxi5911m = reg_1_7&cdxi5180m;
wire cdxi5912m = reg_1_5&cdxi5444m;
wire cdxi5913m = reg_1_3&cdxi5235m;
wire cdxi5914m = reg_1_2&cdxi5127m;
wire cdxi5915m = (cdxi5901m ^ cdxi5902m ^ cdxi5903m ^ cdxi5904m ^ cdxi5905m ^ cdxi5906m ^ cdxi5907m ^ cdxi5908m ^ cdxi5909m ^ cdxi5910m ^ cdxi5911m ^ cdxi5912m ^ cdxi5913m ^ cdxi5914m ^ cdxi5900m);
wire cdxi5916m = reg_1_0&cdxi5915m;
wire cdxi5917m = cdxi5101m&cdxi4790m;
wire cdxi5918m = cdxi4895m&cdxi4753m;
wire cdxi5919m = cdxi4873m&cdxi4850m;
wire cdxi5920m = cdxi4873m&cdxi4851m;
wire cdxi5921m = cdxi5154m&r13m;
wire cdxi5922m = cdxi4934m&r16m;
wire cdxi5923m = cdxi5101m&r17m;
wire cdxi5924m = cdxi5065m&r20m;
wire cdxi5925m = cdxi4895m&r21m;
wire cdxi5926m = cdxi4873m&r27m;
wire cdxi5927m = cdxi4732m&r45m;
wire cdxi5928m = cdxi4742m&r46m;
wire cdxi5929m = cdxi4711m&r52m;
wire cdxi5930m = cdxi4743m&r58m;
wire cdxi5931m = (cdxi88m ^ cdxi5917m ^ cdxi5918m ^ cdxi5919m ^ cdxi5920m ^ cdxi5921m ^ cdxi5922m ^ cdxi5923m ^ cdxi5924m ^ cdxi5925m ^ cdxi5926m ^ cdxi5927m ^ cdxi5928m ^ cdxi5929m ^ cdxi5930m);
wire cdxi5932m = a1&cdxi5931m;
wire cdxi5933m = (reg_1_96);
wire cdxi5934m = reg_1_3&reg_1_6&cdxi4795m;
wire cdxi5935m = reg_1_2&reg_1_6&cdxi4758m;
wire cdxi5936m = reg_1_2&reg_1_3&cdxi4855m;
wire cdxi5937m = reg_1_2&reg_1_3&cdxi4856m;
wire cdxi5938m = reg_1_6&reg_1_7&cdxi4885m;
wire cdxi5939m = reg_1_3&reg_1_7&cdxi4748m;
wire cdxi5940m = reg_1_3&reg_1_6&cdxi4794m;
wire cdxi5941m = reg_1_2&reg_1_7&cdxi4812m;
wire cdxi5942m = reg_1_2&reg_1_6&cdxi4757m;
wire cdxi5943m = reg_1_2&reg_1_3&cdxi4854m;
wire cdxi5944m = reg_1_7&cdxi5197m;
wire cdxi5945m = reg_1_6&cdxi5444m;
wire cdxi5946m = reg_1_3&cdxi5552m;
wire cdxi5947m = reg_1_2&cdxi5692m;
wire cdxi5948m = (cdxi5934m ^ cdxi5935m ^ cdxi5936m ^ cdxi5937m ^ cdxi5938m ^ cdxi5939m ^ cdxi5940m ^ cdxi5941m ^ cdxi5942m ^ cdxi5943m ^ cdxi5944m ^ cdxi5945m ^ cdxi5946m ^ cdxi5947m ^ cdxi5933m);
wire cdxi5949m = reg_1_0&cdxi5948m;
wire cdxi5950m = cdxi4953m&cdxi4742m;
wire cdxi5951m = cdxi4953m&cdxi4744m;
wire cdxi5952m = cdxi5028m&cdxi4817m;
wire cdxi5953m = cdxi5009m&cdxi4772m;
wire cdxi5954m = cdxi5009m&cdxi4773m;
wire cdxi5955m = cdxi4762m&cdxi5050m;
wire cdxi5956m = cdxi4973m&r15m;
wire cdxi5957m = cdxi4953m&r16m;
wire cdxi5958m = cdxi4895m&r22m;
wire cdxi5959m = cdxi5028m&r23m;
wire cdxi5960m = cdxi5009m&r25m;
wire cdxi5961m = cdxi4742m&r47m;
wire cdxi5962m = cdxi4762m&r48m;
wire cdxi5963m = cdxi4722m&r50m;
wire cdxi5964m = cdxi4743m&r59m;
wire cdxi5965m = (cdxi89m ^ cdxi5951m ^ cdxi5952m ^ cdxi5953m ^ cdxi5954m ^ cdxi5955m ^ cdxi5956m ^ cdxi5957m ^ cdxi5958m ^ cdxi5959m ^ cdxi5960m ^ cdxi5961m ^ cdxi5962m ^ cdxi5963m ^ cdxi5964m);
wire cdxi5966m = a1&cdxi5965m;
wire cdxi5967m = (reg_1_97);
wire cdxi5968m = reg_1_4&cdxi5219m;
wire cdxi5969m = reg_1_2&cdxi5146m;
wire cdxi5970m = reg_1_2&cdxi5147m;
wire cdxi5971m = reg_1_2&cdxi5148m;
wire cdxi5972m = reg_1_5&cdxi5059m;
wire cdxi5973m = reg_1_4&cdxi5222m;
wire cdxi5974m = reg_1_4&cdxi5223m;
wire cdxi5975m = reg_1_2&cdxi5149m;
wire cdxi5976m = reg_1_2&cdxi5150m;
wire cdxi5977m = reg_1_2&cdxi5151m;
wire cdxi5978m = reg_1_6&cdxi5038m;
wire cdxi5979m = reg_1_5&cdxi5055m;
wire cdxi5980m = reg_1_4&cdxi5218m;
wire cdxi5981m = reg_1_2&cdxi5145m;
wire cdxi5982m = (cdxi5968m ^ cdxi5969m ^ cdxi5970m ^ cdxi5971m ^ cdxi5972m ^ cdxi5973m ^ cdxi5974m ^ cdxi5975m ^ cdxi5976m ^ cdxi5977m ^ cdxi5978m ^ cdxi5979m ^ cdxi5980m ^ cdxi5981m ^ cdxi5967m);
wire cdxi5983m = reg_1_0&cdxi5982m;
wire cdxi5984m = cdxi4953m&cdxi4790m;
wire cdxi5985m = cdxi5028m&cdxi4839m;
wire cdxi5986m = cdxi5009m&cdxi4781m;
wire cdxi5987m = cdxi5009m&cdxi4782m;
wire cdxi5988m = cdxi4991m&r14m;
wire cdxi5989m = cdxi5064m&r15m;
wire cdxi5990m = cdxi4953m&r17m;
wire cdxi5991m = cdxi5065m&r22m;
wire cdxi5992m = cdxi5028m&r24m;
wire cdxi5993m = cdxi5009m&r26m;
wire cdxi5994m = cdxi4732m&r47m;
wire cdxi5995m = cdxi4762m&r49m;
wire cdxi5996m = cdxi4722m&r51m;
wire cdxi5997m = cdxi4743m&r60m;
wire cdxi5998m = (cdxi90m ^ cdxi5984m ^ cdxi5985m ^ cdxi5986m ^ cdxi5987m ^ cdxi5988m ^ cdxi5989m ^ cdxi5990m ^ cdxi5991m ^ cdxi5992m ^ cdxi5993m ^ cdxi5994m ^ cdxi5995m ^ cdxi5996m ^ cdxi5997m);
wire cdxi5999m = a1&cdxi5998m;
wire cdxi6000m = (reg_1_98);
wire cdxi6001m = reg_1_4&cdxi5236m;
wire cdxi6002m = reg_1_2&cdxi5301m;
wire cdxi6003m = reg_1_2&cdxi5302m;
wire cdxi6004m = reg_1_2&cdxi5303m;
wire cdxi6005m = reg_1_5&cdxi5078m;
wire cdxi6006m = reg_1_4&cdxi5239m;
wire cdxi6007m = reg_1_4&cdxi5240m;
wire cdxi6008m = reg_1_2&cdxi5304m;
wire cdxi6009m = reg_1_2&cdxi5305m;
wire cdxi6010m = reg_1_2&cdxi5306m;
wire cdxi6011m = reg_1_7&cdxi5038m;
wire cdxi6012m = reg_1_5&cdxi5074m;
wire cdxi6013m = reg_1_4&cdxi5235m;
wire cdxi6014m = reg_1_2&cdxi5300m;
wire cdxi6015m = (cdxi6001m ^ cdxi6002m ^ cdxi6003m ^ cdxi6004m ^ cdxi6005m ^ cdxi6006m ^ cdxi6007m ^ cdxi6008m ^ cdxi6009m ^ cdxi6010m ^ cdxi6011m ^ cdxi6012m ^ cdxi6013m ^ cdxi6014m ^ cdxi6000m);
wire cdxi6016m = reg_1_0&cdxi6015m;
wire cdxi6017m = cdxi5136m&cdxi4732m;
wire cdxi6018m = cdxi5136m&cdxi4753m;
wire cdxi6019m = cdxi5101m&cdxi4781m;
wire cdxi6020m = cdxi5083m&cdxi4850m;
wire cdxi6021m = cdxi5083m&cdxi4851m;
wire cdxi6022m = cdxi4742m&cdxi5122m;
wire cdxi6023m = cdxi4991m&r20m;
wire cdxi6024m = cdxi5136m&r21m;
wire cdxi6025m = cdxi4934m&r25m;
wire cdxi6026m = cdxi5101m&r26m;
wire cdxi6027m = cdxi5083m&r27m;
wire cdxi6028m = cdxi4732m&r56m;
wire cdxi6029m = cdxi4742m&r57m;
wire cdxi6030m = cdxi4762m&r58m;
wire cdxi6031m = cdxi4711m&r62m;
wire cdxi6032m = (cdxi96m ^ cdxi6018m ^ cdxi6019m ^ cdxi6020m ^ cdxi6021m ^ cdxi6022m ^ cdxi6023m ^ cdxi6024m ^ cdxi6025m ^ cdxi6026m ^ cdxi6027m ^ cdxi6028m ^ cdxi6029m ^ cdxi6030m ^ cdxi6031m);
wire cdxi6033m = a1&cdxi6032m;
wire cdxi6034m = (reg_1_104);
wire cdxi6035m = reg_1_5&reg_1_6&cdxi4758m;
wire cdxi6036m = reg_1_3&cdxi5164m;
wire cdxi6037m = reg_1_3&cdxi5165m;
wire cdxi6038m = reg_1_3&cdxi5166m;
wire cdxi6039m = reg_1_6&cdxi5131m;
wire cdxi6040m = reg_1_5&reg_1_7&cdxi4812m;
wire cdxi6041m = reg_1_5&reg_1_6&cdxi4757m;
wire cdxi6042m = reg_1_3&cdxi5167m;
wire cdxi6043m = reg_1_3&cdxi5168m;
wire cdxi6044m = reg_1_3&cdxi5169m;
wire cdxi6045m = reg_1_7&cdxi5865m;
wire cdxi6046m = reg_1_6&cdxi5127m;
wire cdxi6047m = reg_1_5&cdxi5692m;
wire cdxi6048m = reg_1_3&cdxi5163m;
wire cdxi6049m = (cdxi6035m ^ cdxi6036m ^ cdxi6037m ^ cdxi6038m ^ cdxi6039m ^ cdxi6040m ^ cdxi6041m ^ cdxi6042m ^ cdxi6043m ^ cdxi6044m ^ cdxi6045m ^ cdxi6046m ^ cdxi6047m ^ cdxi6048m ^ cdxi6034m);
wire cdxi6050m = reg_1_0&cdxi6049m;
wire cdxi6051m = cdxi4915m&cdxi4744m;
wire cdxi6052m = cdxi5009m&cdxi4808m;
wire cdxi6053m = cdxi4873m&cdxi4817m;
wire cdxi6054m = cdxi4873m&cdxi4818m;
wire cdxi6055m = cdxi4973m&r13m;
wire cdxi6056m = cdxi4711m&cdxi5050m;
wire cdxi6057m = cdxi4915m&r16m;
wire cdxi6058m = cdxi4895m&r18m;
wire cdxi6059m = cdxi5009m&r20m;
wire cdxi6060m = cdxi4873m&r23m;
wire cdxi6061m = cdxi4742m&r43m;
wire cdxi6062m = cdxi4722m&r45m;
wire cdxi6063m = cdxi4711m&r48m;
wire cdxi6064m = cdxi4743m&r54m;
wire cdxi6065m = (cdxi84m ^ cdxi6051m ^ cdxi6052m ^ cdxi6053m ^ cdxi6054m ^ cdxi6055m ^ cdxi6056m ^ cdxi6057m ^ cdxi6058m ^ cdxi6059m ^ cdxi6060m ^ cdxi6061m ^ cdxi6062m ^ cdxi6063m ^ cdxi6064m);
wire cdxi6066m = cdxi4712m&cdxi6065m;
wire cdxi6067m = (reg_1_92);
wire cdxi6068m = reg_1_3&cdxi5056m;
wire cdxi6069m = reg_1_2&cdxi5111m;
wire cdxi6070m = reg_1_2&cdxi5112m;
wire cdxi6071m = reg_1_2&cdxi5113m;
wire cdxi6072m = reg_1_4&cdxi5201m;
wire cdxi6073m = reg_1_3&cdxi5059m;
wire cdxi6074m = reg_1_3&cdxi5060m;
wire cdxi6075m = reg_1_2&cdxi5114m;
wire cdxi6076m = reg_1_2&cdxi5115m;
wire cdxi6077m = reg_1_2&cdxi5116m;
wire cdxi6078m = reg_1_6&cdxi5019m;
wire cdxi6079m = reg_1_4&cdxi5197m;
wire cdxi6080m = reg_1_3&cdxi5055m;
wire cdxi6081m = reg_1_2&cdxi5110m;
wire cdxi6082m = (cdxi6068m ^ cdxi6069m ^ cdxi6070m ^ cdxi6071m ^ cdxi6072m ^ cdxi6073m ^ cdxi6074m ^ cdxi6075m ^ cdxi6076m ^ cdxi6077m ^ cdxi6078m ^ cdxi6079m ^ cdxi6080m ^ cdxi6081m ^ cdxi6067m);
wire cdxi6083m = reg_1_1&cdxi6082m;
wire cdxi6084m = cdxi4712m&cdxi5998m;
wire cdxi6085m = reg_1_1&cdxi6015m;
wire cdxi6086m = cdxi4953m&cdxi4753m;
wire cdxi6087m = cdxi5083m&cdxi4839m;
wire cdxi6088m = cdxi4915m&cdxi4781m;
wire cdxi6089m = cdxi4915m&cdxi4782m;
wire cdxi6090m = cdxi4991m&r18m;
wire cdxi6091m = cdxi5064m&r19m;
wire cdxi6092m = cdxi4953m&r21m;
wire cdxi6093m = cdxi4934m&r22m;
wire cdxi6094m = cdxi5083m&r24m;
wire cdxi6095m = cdxi4915m&r26m;
wire cdxi6096m = cdxi4732m&r53m;
wire cdxi6097m = cdxi4762m&r55m;
wire cdxi6098m = cdxi4722m&r57m;
wire cdxi6099m = cdxi4711m&r60m;
wire cdxi6100m = (cdxi94m ^ cdxi6086m ^ cdxi6087m ^ cdxi6088m ^ cdxi6089m ^ cdxi6090m ^ cdxi6091m ^ cdxi6092m ^ cdxi6093m ^ cdxi6094m ^ cdxi6095m ^ cdxi6096m ^ cdxi6097m ^ cdxi6098m ^ cdxi6099m);
wire cdxi6101m = cdxi4712m&cdxi6100m;
wire cdxi6102m = (reg_1_102);
wire cdxi6103m = reg_1_4&cdxi5128m;
wire cdxi6104m = reg_1_3&cdxi5301m;
wire cdxi6105m = reg_1_3&cdxi5302m;
wire cdxi6106m = reg_1_3&cdxi5303m;
wire cdxi6107m = reg_1_5&cdxi5281m;
wire cdxi6108m = reg_1_4&cdxi5131m;
wire cdxi6109m = reg_1_4&cdxi5132m;
wire cdxi6110m = reg_1_3&cdxi5304m;
wire cdxi6111m = reg_1_3&cdxi5305m;
wire cdxi6112m = reg_1_3&cdxi5306m;
wire cdxi6113m = reg_1_7&cdxi5092m;
wire cdxi6114m = reg_1_5&cdxi5277m;
wire cdxi6115m = reg_1_4&cdxi5127m;
wire cdxi6116m = reg_1_3&cdxi5300m;
wire cdxi6117m = (cdxi6103m ^ cdxi6104m ^ cdxi6105m ^ cdxi6106m ^ cdxi6107m ^ cdxi6108m ^ cdxi6109m ^ cdxi6110m ^ cdxi6111m ^ cdxi6112m ^ cdxi6113m ^ cdxi6114m ^ cdxi6115m ^ cdxi6116m ^ cdxi6102m);
wire cdxi6118m = reg_1_1&cdxi6117m;
wire cdxi6119m = cdxi4973m&cdxi4753m;
wire cdxi6120m = cdxi5101m&cdxi4839m;
wire cdxi6121m = cdxi4915m&cdxi4850m;
wire cdxi6122m = cdxi4915m&cdxi4851m;
wire cdxi6123m = cdxi5154m&r18m;
wire cdxi6124m = cdxi5064m&r20m;
wire cdxi6125m = cdxi4973m&r21m;
wire cdxi6126m = cdxi4934m&r23m;
wire cdxi6127m = cdxi5101m&r24m;
wire cdxi6128m = cdxi4915m&r27m;
wire cdxi6129m = cdxi4732m&r54m;
wire cdxi6130m = cdxi4742m&r55m;
wire cdxi6131m = cdxi4722m&r58m;
wire cdxi6132m = cdxi4711m&r61m;
wire cdxi6133m = (cdxi95m ^ cdxi6119m ^ cdxi6120m ^ cdxi6121m ^ cdxi6122m ^ cdxi6123m ^ cdxi6124m ^ cdxi6125m ^ cdxi6126m ^ cdxi6127m ^ cdxi6128m ^ cdxi6129m ^ cdxi6130m ^ cdxi6131m ^ cdxi6132m);
wire cdxi6134m = cdxi4712m&cdxi6133m;
wire cdxi6135m = (reg_1_103);
wire cdxi6136m = reg_1_4&reg_1_6&cdxi4758m;
wire cdxi6137m = reg_1_3&cdxi5259m;
wire cdxi6138m = reg_1_3&cdxi5260m;
wire cdxi6139m = reg_1_3&cdxi5261m;
wire cdxi6140m = reg_1_6&cdxi5281m;
wire cdxi6141m = reg_1_4&reg_1_7&cdxi4812m;
wire cdxi6142m = reg_1_4&reg_1_6&cdxi4757m;
wire cdxi6143m = reg_1_3&cdxi5262m;
wire cdxi6144m = reg_1_3&cdxi5263m;
wire cdxi6145m = reg_1_3&cdxi5264m;
wire cdxi6146m = reg_1_7&cdxi5110m;
wire cdxi6147m = reg_1_6&cdxi5277m;
wire cdxi6148m = reg_1_4&cdxi5692m;
wire cdxi6149m = reg_1_3&cdxi5258m;
wire cdxi6150m = (cdxi6136m ^ cdxi6137m ^ cdxi6138m ^ cdxi6139m ^ cdxi6140m ^ cdxi6141m ^ cdxi6142m ^ cdxi6143m ^ cdxi6144m ^ cdxi6145m ^ cdxi6146m ^ cdxi6147m ^ cdxi6148m ^ cdxi6149m ^ cdxi6135m);
wire cdxi6151m = reg_1_1&cdxi6150m;
wire cdxi6152m = cdxi4953m&cdxi4808m;
wire cdxi6153m = cdxi5083m&cdxi4817m;
wire cdxi6154m = cdxi4915m&cdxi4772m;
wire cdxi6155m = cdxi4915m&cdxi4773m;
wire cdxi6156m = cdxi4762m&cdxi5105m;
wire cdxi6157m = cdxi4973m&r19m;
wire cdxi6158m = cdxi4953m&r20m;
wire cdxi6159m = cdxi5101m&r22m;
wire cdxi6160m = cdxi5083m&r23m;
wire cdxi6161m = cdxi4915m&r25m;
wire cdxi6162m = cdxi4742m&r53m;
wire cdxi6163m = cdxi4762m&r54m;
wire cdxi6164m = cdxi4722m&r56m;
wire cdxi6165m = cdxi4711m&r59m;
wire cdxi6166m = (cdxi93m ^ cdxi6152m ^ cdxi6153m ^ cdxi6154m ^ cdxi6155m ^ cdxi6156m ^ cdxi6157m ^ cdxi6158m ^ cdxi6159m ^ cdxi6160m ^ cdxi6161m ^ cdxi6162m ^ cdxi6163m ^ cdxi6164m ^ cdxi6165m);
wire cdxi6167m = cdxi4743m&cdxi6166m;
wire cdxi6168m = (reg_1_101);
wire cdxi6169m = reg_1_4&reg_1_5&cdxi4813m;
wire cdxi6170m = reg_1_3&cdxi5146m;
wire cdxi6171m = reg_1_3&cdxi5147m;
wire cdxi6172m = reg_1_3&cdxi5148m;
wire cdxi6173m = reg_1_5&cdxi5114m;
wire cdxi6174m = reg_1_4&reg_1_6&cdxi4830m;
wire cdxi6175m = reg_1_4&reg_1_5&cdxi4812m;
wire cdxi6176m = reg_1_3&cdxi5149m;
wire cdxi6177m = reg_1_3&cdxi5150m;
wire cdxi6178m = reg_1_3&cdxi5151m;
wire cdxi6179m = reg_1_6&cdxi5092m;
wire cdxi6180m = reg_1_5&cdxi5110m;
wire cdxi6181m = reg_1_4&cdxi5865m;
wire cdxi6182m = reg_1_3&cdxi5145m;
wire cdxi6183m = (cdxi6169m ^ cdxi6170m ^ cdxi6171m ^ cdxi6172m ^ cdxi6173m ^ cdxi6174m ^ cdxi6175m ^ cdxi6176m ^ cdxi6177m ^ cdxi6178m ^ cdxi6179m ^ cdxi6180m ^ cdxi6181m ^ cdxi6182m ^ cdxi6168m);
wire cdxi6184m = reg_1_2&cdxi6183m;
wire cdxi6185m = cdxi4743m&cdxi6100m;
wire cdxi6186m = reg_1_2&cdxi6117m;
wire cdxi6187m = cdxi4743m&cdxi6133m;
wire cdxi6188m = reg_1_2&cdxi6150m;
wire cdxi6189m = cdxi4743m&cdxi6032m;
wire cdxi6190m = reg_1_2&cdxi6049m;
wire cdxi6191m = cdxi5136m&cdxi4839m;
wire cdxi6192m = cdxi4973m&cdxi4781m;
wire cdxi6193m = cdxi4953m&cdxi4850m;
wire cdxi6194m = cdxi4953m&cdxi4851m;
wire cdxi6195m = cdxi5154m&r22m;
wire cdxi6196m = cdxi4991m&r23m;
wire cdxi6197m = cdxi5136m&r24m;
wire cdxi6198m = cdxi5064m&r25m;
wire cdxi6199m = cdxi4973m&r26m;
wire cdxi6200m = cdxi4953m&r27m;
wire cdxi6201m = cdxi4732m&r59m;
wire cdxi6202m = cdxi4742m&r60m;
wire cdxi6203m = cdxi4762m&r61m;
wire cdxi6204m = cdxi4722m&r62m;
wire cdxi6205m = (cdxi97m ^ cdxi6191m ^ cdxi6192m ^ cdxi6193m ^ cdxi6194m ^ cdxi6195m ^ cdxi6196m ^ cdxi6197m ^ cdxi6198m ^ cdxi6199m ^ cdxi6200m ^ cdxi6201m ^ cdxi6202m ^ cdxi6203m ^ cdxi6204m);
wire cdxi6206m = cdxi4711m&cdxi6205m;
wire cdxi6207m = (reg_1_105);
wire cdxi6208m = reg_1_5&cdxi5259m;
wire cdxi6209m = reg_1_4&cdxi5164m;
wire cdxi6210m = reg_1_4&cdxi5165m;
wire cdxi6211m = reg_1_4&cdxi5166m;
wire cdxi6212m = reg_1_6&cdxi5304m;
wire cdxi6213m = reg_1_5&cdxi5262m;
wire cdxi6214m = reg_1_5&cdxi5263m;
wire cdxi6215m = reg_1_4&cdxi5167m;
wire cdxi6216m = reg_1_4&cdxi5168m;
wire cdxi6217m = reg_1_4&cdxi5169m;
wire cdxi6218m = reg_1_7&cdxi5145m;
wire cdxi6219m = reg_1_6&cdxi5300m;
wire cdxi6220m = reg_1_5&cdxi5258m;
wire cdxi6221m = reg_1_4&cdxi5163m;
wire cdxi6222m = (cdxi6208m ^ cdxi6209m ^ cdxi6210m ^ cdxi6211m ^ cdxi6212m ^ cdxi6213m ^ cdxi6214m ^ cdxi6215m ^ cdxi6216m ^ cdxi6217m ^ cdxi6218m ^ cdxi6219m ^ cdxi6220m ^ cdxi6221m ^ cdxi6207m);
wire cdxi6223m = reg_1_3&cdxi6222m;
wire cdxi6224m = cdxi4873m&cdxi4953m;
wire cdxi6225m = cdxi4874m&cdxi4953m;
wire cdxi6226m = cdxi4875m&cdxi4953m;
wire cdxi6227m = cdxi5314m&cdxi4762m;
wire cdxi6228m = cdxi4712m&cdxi5311m;
wire cdxi6229m = cdxi4873m&cdxi4955m;
wire cdxi6230m = cdxi4874m&cdxi5029m;
wire cdxi6231m = cdxi4875m&cdxi5084m;
wire cdxi6232m = cdxi5314m&cdxi4763m;
wire cdxi6233m = cdxi5314m&cdxi4764m;
wire cdxi6234m = cdxi5779m&r7m;
wire cdxi6235m = cdxi5780m&r8m;
wire cdxi6236m = cdxi4873m&cdxi4958m;
wire cdxi6237m = cdxi4873m&cdxi4959m;
wire cdxi6238m = cdxi4916m&cdxi5175m;
wire cdxi6239m = cdxi4874m&cdxi5032m;
wire cdxi6240m = cdxi4874m&cdxi5033m;
wire cdxi6241m = cdxi4875m&cdxi5087m;
wire cdxi6242m = cdxi4875m&cdxi5088m;
wire cdxi6243m = cdxi5314m&r22m;
wire cdxi6244m = cdxi4953m&r28m;
wire cdxi6245m = cdxi5083m&r29m;
wire cdxi6246m = cdxi4915m&r30m;
wire cdxi6247m = cdxi5028m&r33m;
wire cdxi6248m = cdxi5009m&r34m;
wire cdxi6249m = cdxi4873m&r37m;
wire cdxi6250m = cdxi4954m&r43m;
wire cdxi6251m = cdxi4916m&r44m;
wire cdxi6252m = cdxi4874m&r47m;
wire cdxi6253m = cdxi4875m&r53m;
wire cdxi6254m = cdxi4762m&r63m;
wire cdxi6255m = cdxi4722m&r64m;
wire cdxi6256m = cdxi4711m&r67m;
wire cdxi6257m = cdxi4743m&r73m;
wire cdxi6258m = cdxi4712m&r83m;
wire cdxi6259m = (cdxi98m ^ cdxi6229m ^ cdxi6230m ^ cdxi6231m ^ cdxi6232m ^ cdxi6233m ^ cdxi6234m ^ cdxi6235m ^ cdxi6236m ^ cdxi6237m ^ cdxi6238m ^ cdxi6239m ^ cdxi6240m ^ cdxi6241m ^ cdxi6242m ^ cdxi6243m ^ cdxi6244m ^ cdxi6245m ^ cdxi6246m ^ cdxi6247m ^ cdxi6248m ^ cdxi6249m ^ cdxi6250m ^ cdxi6251m ^ cdxi6252m ^ cdxi6253m ^ cdxi6254m ^ cdxi6255m ^ cdxi6256m ^ cdxi6257m ^ cdxi6258m);
wire cdxi6260m = a1&cdxi6259m;
wire cdxi6261m = (reg_1_75);
wire cdxi6262m = (reg_1_81);
wire cdxi6263m = (reg_1_106);
wire cdxi6264m = reg_1_2&reg_1_3&cdxi4965m;
wire cdxi6265m = reg_1_1&cdxi5798m;
wire cdxi6266m = reg_1_1&cdxi5799m;
wire cdxi6267m = reg_1_1&cdxi5800m;
wire cdxi6268m = reg_1_1&cdxi5801m;
wire cdxi6269m = reg_1_3&reg_1_4&reg_1_5&cdxi4884m;
wire cdxi6270m = reg_1_2&reg_1_4&reg_1_5&cdxi4717m;
wire cdxi6271m = reg_1_2&reg_1_3&cdxi4968m;
wire cdxi6272m = reg_1_2&reg_1_3&cdxi4969m;
wire cdxi6273m = reg_1_1&cdxi5802m;
wire cdxi6274m = reg_1_1&cdxi5803m;
wire cdxi6275m = reg_1_1&cdxi5804m;
wire cdxi6276m = reg_1_1&cdxi5805m;
wire cdxi6277m = reg_1_1&cdxi5806m;
wire cdxi6278m = reg_1_1&cdxi5807m;
wire cdxi6279m = reg_1_4&cdxi5381m;
wire cdxi6280m = reg_1_3&reg_1_5&cdxi5331m;
wire cdxi6281m = reg_1_3&reg_1_4&cdxi5368m;
wire cdxi6282m = reg_1_2&reg_1_5&cdxi4925m;
wire cdxi6283m = reg_1_2&reg_1_4&cdxi5369m;
wire cdxi6284m = reg_1_2&reg_1_3&cdxi4964m;
wire cdxi6285m = reg_1_1&cdxi5808m;
wire cdxi6286m = reg_1_1&cdxi5809m;
wire cdxi6287m = reg_1_1&cdxi5810m;
wire cdxi6288m = reg_1_1&cdxi5811m;
wire cdxi6289m = reg_1_5&cdxi5332m;
wire cdxi6290m = reg_1_4&cdxi5370m;
wire cdxi6291m = reg_1_3&cdxi6261m;
wire cdxi6292m = reg_1_2&cdxi6262m;
wire cdxi6293m = reg_1_1&cdxi5797m;
wire cdxi6294m = (cdxi6264m ^ cdxi6265m ^ cdxi6266m ^ cdxi6267m ^ cdxi6268m ^ cdxi6269m ^ cdxi6270m ^ cdxi6271m ^ cdxi6272m ^ cdxi6273m ^ cdxi6274m ^ cdxi6275m ^ cdxi6276m ^ cdxi6277m ^ cdxi6278m ^ cdxi6279m ^ cdxi6280m ^ cdxi6281m ^ cdxi6282m ^ cdxi6283m ^ cdxi6284m ^ cdxi6285m ^ cdxi6286m ^ cdxi6287m ^ cdxi6288m ^ cdxi6289m ^ cdxi6290m ^ cdxi6291m ^ cdxi6292m ^ cdxi6293m ^ cdxi6263m);
wire cdxi6295m = reg_1_0&cdxi6294m;
wire cdxi6296m = cdxi4873m&cdxi4973m;
wire cdxi6297m = cdxi4874m&cdxi4973m;
wire cdxi6298m = cdxi4875m&cdxi4973m;
wire cdxi6299m = cdxi5314m&cdxi4742m;
wire cdxi6300m = cdxi4873m&cdxi4974m;
wire cdxi6301m = cdxi4874m&cdxi5047m;
wire cdxi6302m = cdxi4875m&cdxi5102m;
wire cdxi6303m = cdxi5314m&cdxi4817m;
wire cdxi6304m = cdxi5314m&cdxi4818m;
wire cdxi6305m = cdxi4915m&cdxi4900m;
wire cdxi6306m = cdxi5462m&r8m;
wire cdxi6307m = cdxi4873m&cdxi4977m;
wire cdxi6308m = cdxi4873m&cdxi4978m;
wire cdxi6309m = cdxi4916m&cdxi5192m;
wire cdxi6310m = cdxi4874m&cdxi5050m;
wire cdxi6311m = cdxi4874m&cdxi5051m;
wire cdxi6312m = cdxi4875m&cdxi5105m;
wire cdxi6313m = cdxi4875m&cdxi5106m;
wire cdxi6314m = cdxi5314m&r23m;
wire cdxi6315m = cdxi4973m&r28m;
wire cdxi6316m = cdxi5101m&r29m;
wire cdxi6317m = cdxi4915m&r31m;
wire cdxi6318m = cdxi4895m&r33m;
wire cdxi6319m = cdxi5009m&r35m;
wire cdxi6320m = cdxi4873m&r38m;
wire cdxi6321m = cdxi4896m&r43m;
wire cdxi6322m = cdxi4916m&r45m;
wire cdxi6323m = cdxi4874m&r48m;
wire cdxi6324m = cdxi4875m&r54m;
wire cdxi6325m = cdxi4742m&r63m;
wire cdxi6326m = cdxi4722m&r65m;
wire cdxi6327m = cdxi4711m&r68m;
wire cdxi6328m = cdxi4743m&r74m;
wire cdxi6329m = cdxi4712m&r84m;
wire cdxi6330m = (cdxi99m ^ cdxi6300m ^ cdxi6301m ^ cdxi6302m ^ cdxi6303m ^ cdxi6304m ^ cdxi6305m ^ cdxi6306m ^ cdxi6307m ^ cdxi6308m ^ cdxi6309m ^ cdxi6310m ^ cdxi6311m ^ cdxi6312m ^ cdxi6313m ^ cdxi6314m ^ cdxi6315m ^ cdxi6316m ^ cdxi6317m ^ cdxi6318m ^ cdxi6319m ^ cdxi6320m ^ cdxi6321m ^ cdxi6322m ^ cdxi6323m ^ cdxi6324m ^ cdxi6325m ^ cdxi6326m ^ cdxi6327m ^ cdxi6328m ^ cdxi6329m);
wire cdxi6331m = a1&cdxi6330m;
wire cdxi6332m = (reg_1_107);
wire cdxi6333m = reg_1_2&cdxi5588m;
wire cdxi6334m = reg_1_1&cdxi6068m;
wire cdxi6335m = reg_1_1&cdxi6069m;
wire cdxi6336m = reg_1_1&cdxi6070m;
wire cdxi6337m = reg_1_1&cdxi6071m;
wire cdxi6338m = reg_1_3&cdxi5485m;
wire cdxi6339m = reg_1_2&cdxi5592m;
wire cdxi6340m = reg_1_2&cdxi5593m;
wire cdxi6341m = reg_1_2&cdxi5594m;
wire cdxi6342m = reg_1_1&cdxi6072m;
wire cdxi6343m = reg_1_1&cdxi6073m;
wire cdxi6344m = reg_1_1&cdxi6074m;
wire cdxi6345m = reg_1_1&cdxi6075m;
wire cdxi6346m = reg_1_1&cdxi6076m;
wire cdxi6347m = reg_1_1&cdxi6077m;
wire cdxi6348m = reg_1_4&cdxi5418m;
wire cdxi6349m = reg_1_3&cdxi5491m;
wire cdxi6350m = reg_1_3&cdxi5492m;
wire cdxi6351m = reg_1_2&cdxi5598m;
wire cdxi6352m = reg_1_2&cdxi5599m;
wire cdxi6353m = reg_1_2&cdxi5600m;
wire cdxi6354m = reg_1_1&cdxi6078m;
wire cdxi6355m = reg_1_1&cdxi6079m;
wire cdxi6356m = reg_1_1&cdxi6080m;
wire cdxi6357m = reg_1_1&cdxi6081m;
wire cdxi6358m = reg_1_6&cdxi5332m;
wire cdxi6359m = reg_1_4&cdxi5407m;
wire cdxi6360m = reg_1_3&cdxi5480m;
wire cdxi6361m = reg_1_2&cdxi5587m;
wire cdxi6362m = reg_1_1&cdxi6067m;
wire cdxi6363m = (cdxi6333m ^ cdxi6334m ^ cdxi6335m ^ cdxi6336m ^ cdxi6337m ^ cdxi6338m ^ cdxi6339m ^ cdxi6340m ^ cdxi6341m ^ cdxi6342m ^ cdxi6343m ^ cdxi6344m ^ cdxi6345m ^ cdxi6346m ^ cdxi6347m ^ cdxi6348m ^ cdxi6349m ^ cdxi6350m ^ cdxi6351m ^ cdxi6352m ^ cdxi6353m ^ cdxi6354m ^ cdxi6355m ^ cdxi6356m ^ cdxi6357m ^ cdxi6358m ^ cdxi6359m ^ cdxi6360m ^ cdxi6361m ^ cdxi6362m ^ cdxi6332m);
wire cdxi6364m = reg_1_0&cdxi6363m;
wire cdxi6365m = cdxi4873m&cdxi5136m;
wire cdxi6366m = cdxi4874m&cdxi5136m;
wire cdxi6367m = cdxi4875m&cdxi5136m;
wire cdxi6368m = cdxi6365m&r0m;
wire cdxi6369m = cdxi4874m&cdxi5210m;
wire cdxi6370m = cdxi5351m&cdxi4808m;
wire cdxi6371m = cdxi5314m&cdxi4772m;
wire cdxi6372m = cdxi5314m&cdxi4773m;
wire cdxi6373m = cdxi5083m&cdxi4900m;
wire cdxi6374m = cdxi5497m&r8m;
wire cdxi6375m = cdxi5387m&r10m;
wire cdxi6376m = cdxi5349m&r11m;
wire cdxi6377m = cdxi4954m&cdxi5192m;
wire cdxi6378m = cdxi4874m&cdxi5213m;
wire cdxi6379m = cdxi4874m&cdxi5214m;
wire cdxi6380m = cdxi5389m&r19m;
wire cdxi6381m = cdxi5351m&r20m;
wire cdxi6382m = cdxi5314m&r25m;
wire cdxi6383m = cdxi5136m&r28m;
wire cdxi6384m = cdxi5101m&r30m;
wire cdxi6385m = cdxi5083m&r31m;
wire cdxi6386m = cdxi4895m&r34m;
wire cdxi6387m = cdxi5028m&r35m;
wire cdxi6388m = cdxi4873m&r40m;
wire cdxi6389m = cdxi4896m&r44m;
wire cdxi6390m = cdxi4954m&r45m;
wire cdxi6391m = cdxi4874m&r50m;
wire cdxi6392m = cdxi4875m&r56m;
wire cdxi6393m = cdxi4742m&r64m;
wire cdxi6394m = cdxi4762m&r65m;
wire cdxi6395m = cdxi4711m&r70m;
wire cdxi6396m = cdxi4743m&r76m;
wire cdxi6397m = cdxi4712m&r86m;
wire cdxi6398m = (cdxi101m ^ cdxi6368m ^ cdxi6369m ^ cdxi6370m ^ cdxi6371m ^ cdxi6372m ^ cdxi6373m ^ cdxi6374m ^ cdxi6375m ^ cdxi6376m ^ cdxi6377m ^ cdxi6378m ^ cdxi6379m ^ cdxi6380m ^ cdxi6381m ^ cdxi6382m ^ cdxi6383m ^ cdxi6384m ^ cdxi6385m ^ cdxi6386m ^ cdxi6387m ^ cdxi6388m ^ cdxi6389m ^ cdxi6390m ^ cdxi6391m ^ cdxi6392m ^ cdxi6393m ^ cdxi6394m ^ cdxi6395m ^ cdxi6396m ^ cdxi6397m);
wire cdxi6399m = a1&cdxi6398m;
wire cdxi6400m = (reg_1_84);
wire cdxi6401m = (reg_1_109);
wire cdxi6402m = reg_1_2&reg_1_3&reg_1_5&reg_1_6&cdxi4664m;
wire cdxi6403m = reg_1_1&cdxi5867m;
wire cdxi6404m = reg_1_1&cdxi5868m;
wire cdxi6405m = reg_1_1&cdxi5869m;
wire cdxi6406m = reg_1_1&cdxi5870m;
wire cdxi6407m = reg_1_3&cdxi5521m;
wire cdxi6408m = reg_1_2&reg_1_5&reg_1_6&cdxi4717m;
wire cdxi6409m = reg_1_2&reg_1_3&reg_1_6&cdxi4963m;
wire cdxi6410m = reg_1_2&reg_1_3&reg_1_5&cdxi4905m;
wire cdxi6411m = reg_1_1&cdxi5871m;
wire cdxi6412m = reg_1_1&cdxi5872m;
wire cdxi6413m = reg_1_1&cdxi5873m;
wire cdxi6414m = reg_1_1&cdxi5874m;
wire cdxi6415m = reg_1_1&cdxi5875m;
wire cdxi6416m = reg_1_1&cdxi5876m;
wire cdxi6417m = reg_1_5&cdxi5418m;
wire cdxi6418m = reg_1_3&cdxi5527m;
wire cdxi6419m = reg_1_3&cdxi5528m;
wire cdxi6420m = reg_1_2&reg_1_6&cdxi5369m;
wire cdxi6421m = reg_1_2&reg_1_5&cdxi5406m;
wire cdxi6422m = reg_1_2&reg_1_3&cdxi5515m;
wire cdxi6423m = reg_1_1&cdxi5877m;
wire cdxi6424m = reg_1_1&cdxi5878m;
wire cdxi6425m = reg_1_1&cdxi5879m;
wire cdxi6426m = reg_1_1&cdxi5880m;
wire cdxi6427m = reg_1_6&cdxi5370m;
wire cdxi6428m = reg_1_5&cdxi5407m;
wire cdxi6429m = reg_1_3&cdxi5516m;
wire cdxi6430m = reg_1_2&cdxi6400m;
wire cdxi6431m = reg_1_1&cdxi5866m;
wire cdxi6432m = (cdxi6402m ^ cdxi6403m ^ cdxi6404m ^ cdxi6405m ^ cdxi6406m ^ cdxi6407m ^ cdxi6408m ^ cdxi6409m ^ cdxi6410m ^ cdxi6411m ^ cdxi6412m ^ cdxi6413m ^ cdxi6414m ^ cdxi6415m ^ cdxi6416m ^ cdxi6417m ^ cdxi6418m ^ cdxi6419m ^ cdxi6420m ^ cdxi6421m ^ cdxi6422m ^ cdxi6423m ^ cdxi6424m ^ cdxi6425m ^ cdxi6426m ^ cdxi6427m ^ cdxi6428m ^ cdxi6429m ^ cdxi6430m ^ cdxi6431m ^ cdxi6401m);
wire cdxi6433m = reg_1_0&cdxi6432m;
wire cdxi6434m = cdxi4873m&cdxi4991m;
wire cdxi6435m = cdxi4874m&cdxi4991m;
wire cdxi6436m = cdxi4875m&cdxi4991m;
wire cdxi6437m = cdxi5314m&cdxi4732m;
wire cdxi6438m = cdxi4873m&cdxi4992m;
wire cdxi6439m = cdxi4874m&cdxi5227m;
wire cdxi6440m = cdxi4875m&cdxi5119m;
wire cdxi6441m = cdxi5314m&cdxi4781m;
wire cdxi6442m = cdxi5314m&cdxi4782m;
wire cdxi6443m = cdxi5640m&r7m;
wire cdxi6444m = cdxi5028m&cdxi4939m;
wire cdxi6445m = cdxi4873m&cdxi4995m;
wire cdxi6446m = cdxi4873m&cdxi4996m;
wire cdxi6447m = cdxi5641m&r13m;
wire cdxi6448m = cdxi4874m&cdxi5230m;
wire cdxi6449m = cdxi4874m&cdxi5231m;
wire cdxi6450m = cdxi4875m&cdxi5122m;
wire cdxi6451m = cdxi4875m&cdxi5123m;
wire cdxi6452m = cdxi5314m&r26m;
wire cdxi6453m = cdxi4991m&r28m;
wire cdxi6454m = cdxi4934m&r30m;
wire cdxi6455m = cdxi5083m&r32m;
wire cdxi6456m = cdxi5065m&r34m;
wire cdxi6457m = cdxi5028m&r36m;
wire cdxi6458m = cdxi4873m&r41m;
wire cdxi6459m = cdxi4935m&r44m;
wire cdxi6460m = cdxi4954m&r46m;
wire cdxi6461m = cdxi4874m&r51m;
wire cdxi6462m = cdxi4875m&r57m;
wire cdxi6463m = cdxi4732m&r64m;
wire cdxi6464m = cdxi4762m&r66m;
wire cdxi6465m = cdxi4711m&r71m;
wire cdxi6466m = cdxi4743m&r77m;
wire cdxi6467m = cdxi4712m&r87m;
wire cdxi6468m = (cdxi102m ^ cdxi6438m ^ cdxi6439m ^ cdxi6440m ^ cdxi6441m ^ cdxi6442m ^ cdxi6443m ^ cdxi6444m ^ cdxi6445m ^ cdxi6446m ^ cdxi6447m ^ cdxi6448m ^ cdxi6449m ^ cdxi6450m ^ cdxi6451m ^ cdxi6452m ^ cdxi6453m ^ cdxi6454m ^ cdxi6455m ^ cdxi6456m ^ cdxi6457m ^ cdxi6458m ^ cdxi6459m ^ cdxi6460m ^ cdxi6461m ^ cdxi6462m ^ cdxi6463m ^ cdxi6464m ^ cdxi6465m ^ cdxi6466m ^ cdxi6467m);
wire cdxi6469m = a1&cdxi6468m;
wire cdxi6470m = (reg_1_79);
wire cdxi6471m = (reg_1_110);
wire cdxi6472m = reg_1_2&cdxi5659m;
wire cdxi6473m = reg_1_1&cdxi5901m;
wire cdxi6474m = reg_1_1&cdxi5902m;
wire cdxi6475m = reg_1_1&cdxi5903m;
wire cdxi6476m = reg_1_1&cdxi5904m;
wire cdxi6477m = reg_1_3&reg_1_5&reg_1_7&cdxi4884m;
wire cdxi6478m = reg_1_2&cdxi5663m;
wire cdxi6479m = reg_1_2&cdxi5664m;
wire cdxi6480m = reg_1_2&cdxi5665m;
wire cdxi6481m = reg_1_1&cdxi5905m;
wire cdxi6482m = reg_1_1&cdxi5906m;
wire cdxi6483m = reg_1_1&cdxi5907m;
wire cdxi6484m = reg_1_1&cdxi5908m;
wire cdxi6485m = reg_1_1&cdxi5909m;
wire cdxi6486m = reg_1_1&cdxi5910m;
wire cdxi6487m = reg_1_5&cdxi5456m;
wire cdxi6488m = reg_1_3&reg_1_7&cdxi5368m;
wire cdxi6489m = reg_1_3&reg_1_5&cdxi5443m;
wire cdxi6490m = reg_1_2&cdxi5669m;
wire cdxi6491m = reg_1_2&cdxi5670m;
wire cdxi6492m = reg_1_2&cdxi5671m;
wire cdxi6493m = reg_1_1&cdxi5911m;
wire cdxi6494m = reg_1_1&cdxi5912m;
wire cdxi6495m = reg_1_1&cdxi5913m;
wire cdxi6496m = reg_1_1&cdxi5914m;
wire cdxi6497m = reg_1_7&cdxi5370m;
wire cdxi6498m = reg_1_5&cdxi5445m;
wire cdxi6499m = reg_1_3&cdxi6470m;
wire cdxi6500m = reg_1_2&cdxi5658m;
wire cdxi6501m = reg_1_1&cdxi5900m;
wire cdxi6502m = (cdxi6472m ^ cdxi6473m ^ cdxi6474m ^ cdxi6475m ^ cdxi6476m ^ cdxi6477m ^ cdxi6478m ^ cdxi6479m ^ cdxi6480m ^ cdxi6481m ^ cdxi6482m ^ cdxi6483m ^ cdxi6484m ^ cdxi6485m ^ cdxi6486m ^ cdxi6487m ^ cdxi6488m ^ cdxi6489m ^ cdxi6490m ^ cdxi6491m ^ cdxi6492m ^ cdxi6493m ^ cdxi6494m ^ cdxi6495m ^ cdxi6496m ^ cdxi6497m ^ cdxi6498m ^ cdxi6499m ^ cdxi6500m ^ cdxi6501m ^ cdxi6471m);
wire cdxi6503m = reg_1_0&cdxi6502m;
wire cdxi6504m = cdxi5780m&cdxi4742m;
wire cdxi6505m = cdxi4916m&cdxi5136m;
wire cdxi6506m = cdxi6504m&r0m;
wire cdxi6507m = cdxi4916m&cdxi5210m;
wire cdxi6508m = cdxi4875m&cdxi5137m;
wire cdxi6509m = cdxi4875m&cdxi5138m;
wire cdxi6510m = cdxi4875m&cdxi5139m;
wire cdxi6511m = cdxi4953m&cdxi4900m;
wire cdxi6512m = cdxi5028m&cdxi4977m;
wire cdxi6513m = cdxi5462m&r10m;
wire cdxi6514m = cdxi5780m&r11m;
wire cdxi6515m = cdxi4954m&cdxi5050m;
wire cdxi6516m = cdxi4916m&cdxi5213m;
wire cdxi6517m = cdxi4916m&cdxi5214m;
wire cdxi6518m = cdxi4875m&cdxi5140m;
wire cdxi6519m = cdxi4875m&cdxi5141m;
wire cdxi6520m = cdxi4875m&cdxi5142m;
wire cdxi6521m = cdxi5136m&r29m;
wire cdxi6522m = cdxi4973m&r30m;
wire cdxi6523m = cdxi4953m&r31m;
wire cdxi6524m = cdxi4895m&r37m;
wire cdxi6525m = cdxi5028m&r38m;
wire cdxi6526m = cdxi5009m&r40m;
wire cdxi6527m = cdxi4896m&r47m;
wire cdxi6528m = cdxi4954m&r48m;
wire cdxi6529m = cdxi4916m&r50m;
wire cdxi6530m = cdxi4875m&r59m;
wire cdxi6531m = cdxi4742m&r67m;
wire cdxi6532m = cdxi4762m&r68m;
wire cdxi6533m = cdxi4722m&r70m;
wire cdxi6534m = cdxi4743m&r79m;
wire cdxi6535m = cdxi4712m&r89m;
wire cdxi6536m = (cdxi104m ^ cdxi6506m ^ cdxi6507m ^ cdxi6508m ^ cdxi6509m ^ cdxi6510m ^ cdxi6511m ^ cdxi6512m ^ cdxi6513m ^ cdxi6514m ^ cdxi6515m ^ cdxi6516m ^ cdxi6517m ^ cdxi6518m ^ cdxi6519m ^ cdxi6520m ^ cdxi6521m ^ cdxi6522m ^ cdxi6523m ^ cdxi6524m ^ cdxi6525m ^ cdxi6526m ^ cdxi6527m ^ cdxi6528m ^ cdxi6529m ^ cdxi6530m ^ cdxi6531m ^ cdxi6532m ^ cdxi6533m ^ cdxi6534m ^ cdxi6535m);
wire cdxi6537m = a1&cdxi6536m;
wire cdxi6538m = (reg_1_87);
wire cdxi6539m = (reg_1_112);
wire cdxi6540m = reg_1_2&reg_1_4&reg_1_5&reg_1_6&cdxi4664m;
wire cdxi6541m = reg_1_1&cdxi5968m;
wire cdxi6542m = reg_1_1&cdxi5969m;
wire cdxi6543m = reg_1_1&cdxi5970m;
wire cdxi6544m = reg_1_1&cdxi5971m;
wire cdxi6545m = reg_1_4&cdxi5521m;
wire cdxi6546m = reg_1_2&reg_1_5&cdxi4986m;
wire cdxi6547m = reg_1_2&reg_1_4&reg_1_6&cdxi4963m;
wire cdxi6548m = reg_1_2&reg_1_4&reg_1_5&cdxi4905m;
wire cdxi6549m = reg_1_1&cdxi5972m;
wire cdxi6550m = reg_1_1&cdxi5973m;
wire cdxi6551m = reg_1_1&cdxi5974m;
wire cdxi6552m = reg_1_1&cdxi5975m;
wire cdxi6553m = reg_1_1&cdxi5976m;
wire cdxi6554m = reg_1_1&cdxi5977m;
wire cdxi6555m = reg_1_5&cdxi5491m;
wire cdxi6556m = reg_1_4&cdxi5527m;
wire cdxi6557m = reg_1_4&cdxi5528m;
wire cdxi6558m = reg_1_2&reg_1_6&cdxi4964m;
wire cdxi6559m = reg_1_2&reg_1_5&cdxi4982m;
wire cdxi6560m = reg_1_2&reg_1_4&cdxi5515m;
wire cdxi6561m = reg_1_1&cdxi5978m;
wire cdxi6562m = reg_1_1&cdxi5979m;
wire cdxi6563m = reg_1_1&cdxi5980m;
wire cdxi6564m = reg_1_1&cdxi5981m;
wire cdxi6565m = reg_1_6&cdxi6261m;
wire cdxi6566m = reg_1_5&cdxi5480m;
wire cdxi6567m = reg_1_4&cdxi5516m;
wire cdxi6568m = reg_1_2&cdxi6538m;
wire cdxi6569m = reg_1_1&cdxi5967m;
wire cdxi6570m = (cdxi6540m ^ cdxi6541m ^ cdxi6542m ^ cdxi6543m ^ cdxi6544m ^ cdxi6545m ^ cdxi6546m ^ cdxi6547m ^ cdxi6548m ^ cdxi6549m ^ cdxi6550m ^ cdxi6551m ^ cdxi6552m ^ cdxi6553m ^ cdxi6554m ^ cdxi6555m ^ cdxi6556m ^ cdxi6557m ^ cdxi6558m ^ cdxi6559m ^ cdxi6560m ^ cdxi6561m ^ cdxi6562m ^ cdxi6563m ^ cdxi6564m ^ cdxi6565m ^ cdxi6566m ^ cdxi6567m ^ cdxi6568m ^ cdxi6569m ^ cdxi6539m);
wire cdxi6571m = reg_1_0&cdxi6570m;
wire cdxi6572m = cdxi5462m&cdxi4732m;
wire cdxi6573m = cdxi4916m&cdxi5154m;
wire cdxi6574m = cdxi4875m&cdxi5154m;
wire cdxi6575m = cdxi4875m&cdxi5064m;
wire cdxi6576m = cdxi5462m&cdxi4733m;
wire cdxi6577m = cdxi5463m&cdxi4790m;
wire cdxi6578m = cdxi4875m&cdxi5250m;
wire cdxi6579m = cdxi4875m&cdxi5251m;
wire cdxi6580m = cdxi4875m&cdxi5252m;
wire cdxi6581m = cdxi5745m&r7m;
wire cdxi6582m = cdxi5533m&r9m;
wire cdxi6583m = cdxi5814m&r11m;
wire cdxi6584m = cdxi5462m&r12m;
wire cdxi6585m = cdxi4896m&cdxi5069m;
wire cdxi6586m = cdxi5605m&r16m;
wire cdxi6587m = cdxi5463m&r17m;
wire cdxi6588m = cdxi4875m&cdxi5253m;
wire cdxi6589m = cdxi4875m&cdxi5254m;
wire cdxi6590m = cdxi4875m&cdxi5255m;
wire cdxi6591m = cdxi5154m&r29m;
wire cdxi6592m = cdxi5064m&r31m;
wire cdxi6593m = cdxi4973m&r32m;
wire cdxi6594m = cdxi5065m&r38m;
wire cdxi6595m = cdxi4895m&r39m;
wire cdxi6596m = cdxi5009m&r42m;
wire cdxi6597m = cdxi4935m&r48m;
wire cdxi6598m = cdxi4896m&r49m;
wire cdxi6599m = cdxi4916m&r52m;
wire cdxi6600m = cdxi4875m&r61m;
wire cdxi6601m = cdxi4732m&r68m;
wire cdxi6602m = cdxi4742m&r69m;
wire cdxi6603m = cdxi4722m&r72m;
wire cdxi6604m = cdxi4743m&r81m;
wire cdxi6605m = cdxi4712m&r91m;
wire cdxi6606m = (cdxi106m ^ cdxi6576m ^ cdxi6577m ^ cdxi6578m ^ cdxi6579m ^ cdxi6580m ^ cdxi6581m ^ cdxi6582m ^ cdxi6583m ^ cdxi6584m ^ cdxi6585m ^ cdxi6586m ^ cdxi6587m ^ cdxi6588m ^ cdxi6589m ^ cdxi6590m ^ cdxi6591m ^ cdxi6592m ^ cdxi6593m ^ cdxi6594m ^ cdxi6595m ^ cdxi6596m ^ cdxi6597m ^ cdxi6598m ^ cdxi6599m ^ cdxi6600m ^ cdxi6601m ^ cdxi6602m ^ cdxi6603m ^ cdxi6604m ^ cdxi6605m);
wire cdxi6607m = a1&cdxi6606m;
wire cdxi6608m = (reg_1_77);
wire cdxi6609m = (reg_1_99);
wire cdxi6610m = (reg_1_114);
wire cdxi6611m = reg_1_2&cdxi5763m;
wire cdxi6612m = reg_1_1&reg_1_4&reg_1_6&cdxi4795m;
wire cdxi6613m = reg_1_1&reg_1_2&cdxi5259m;
wire cdxi6614m = reg_1_1&reg_1_2&cdxi5260m;
wire cdxi6615m = reg_1_1&reg_1_2&cdxi5261m;
wire cdxi6616m = reg_1_4&cdxi5558m;
wire cdxi6617m = reg_1_2&cdxi5767m;
wire cdxi6618m = reg_1_2&cdxi5768m;
wire cdxi6619m = reg_1_2&cdxi5769m;
wire cdxi6620m = reg_1_1&reg_1_6&cdxi5078m;
wire cdxi6621m = reg_1_1&reg_1_4&reg_1_7&cdxi4748m;
wire cdxi6622m = reg_1_1&reg_1_4&reg_1_6&cdxi4794m;
wire cdxi6623m = reg_1_1&reg_1_2&cdxi5262m;
wire cdxi6624m = reg_1_1&reg_1_2&cdxi5263m;
wire cdxi6625m = reg_1_1&reg_1_2&cdxi5264m;
wire cdxi6626m = reg_1_6&reg_1_7&cdxi5331m;
wire cdxi6627m = reg_1_4&cdxi5564m;
wire cdxi6628m = reg_1_4&cdxi5565m;
wire cdxi6629m = reg_1_2&cdxi5773m;
wire cdxi6630m = reg_1_2&cdxi5774m;
wire cdxi6631m = reg_1_2&cdxi5775m;
wire cdxi6632m = reg_1_1&reg_1_7&cdxi5055m;
wire cdxi6633m = reg_1_1&reg_1_6&cdxi5074m;
wire cdxi6634m = reg_1_1&reg_1_4&cdxi5552m;
wire cdxi6635m = reg_1_1&reg_1_2&cdxi5258m;
wire cdxi6636m = reg_1_7&cdxi5480m;
wire cdxi6637m = reg_1_6&cdxi6608m;
wire cdxi6638m = reg_1_4&cdxi5553m;
wire cdxi6639m = reg_1_2&cdxi5762m;
wire cdxi6640m = reg_1_1&cdxi6609m;
wire cdxi6641m = (cdxi6611m ^ cdxi6612m ^ cdxi6613m ^ cdxi6614m ^ cdxi6615m ^ cdxi6616m ^ cdxi6617m ^ cdxi6618m ^ cdxi6619m ^ cdxi6620m ^ cdxi6621m ^ cdxi6622m ^ cdxi6623m ^ cdxi6624m ^ cdxi6625m ^ cdxi6626m ^ cdxi6627m ^ cdxi6628m ^ cdxi6629m ^ cdxi6630m ^ cdxi6631m ^ cdxi6632m ^ cdxi6633m ^ cdxi6634m ^ cdxi6635m ^ cdxi6636m ^ cdxi6637m ^ cdxi6638m ^ cdxi6639m ^ cdxi6640m ^ cdxi6610m);
wire cdxi6642m = reg_1_0&cdxi6641m;
wire cdxi6643m = cdxi5028m&cdxi5154m;
wire cdxi6644m = cdxi4954m&cdxi5154m;
wire cdxi6645m = cdxi5497m&cdxi4733m;
wire cdxi6646m = cdxi5498m&cdxi4790m;
wire cdxi6647m = cdxi4875m&cdxi5155m;
wire cdxi6648m = cdxi4875m&cdxi5156m;
wire cdxi6649m = cdxi4875m&cdxi5157m;
wire cdxi6650m = cdxi6017m&r7m;
wire cdxi6651m = cdxi4895m&cdxi4995m;
wire cdxi6652m = cdxi5883m&r11m;
wire cdxi6653m = cdxi5497m&r12m;
wire cdxi6654m = cdxi4896m&cdxi5230m;
wire cdxi6655m = cdxi5641m&r16m;
wire cdxi6656m = cdxi5498m&r17m;
wire cdxi6657m = cdxi4875m&cdxi5158m;
wire cdxi6658m = cdxi4875m&cdxi5159m;
wire cdxi6659m = cdxi4875m&cdxi5160m;
wire cdxi6660m = cdxi5154m&r30m;
wire cdxi6661m = cdxi4991m&r31m;
wire cdxi6662m = cdxi5136m&r32m;
wire cdxi6663m = cdxi5065m&r40m;
wire cdxi6664m = cdxi4895m&r41m;
wire cdxi6665m = cdxi5028m&r42m;
wire cdxi6666m = cdxi4935m&r50m;
wire cdxi6667m = cdxi4896m&r51m;
wire cdxi6668m = cdxi4954m&r52m;
wire cdxi6669m = cdxi4875m&r62m;
wire cdxi6670m = cdxi4732m&r70m;
wire cdxi6671m = cdxi4742m&r71m;
wire cdxi6672m = cdxi4762m&r72m;
wire cdxi6673m = cdxi4743m&r82m;
wire cdxi6674m = cdxi4712m&r92m;
wire cdxi6675m = (cdxi107m ^ cdxi6645m ^ cdxi6646m ^ cdxi6647m ^ cdxi6648m ^ cdxi6649m ^ cdxi6650m ^ cdxi6651m ^ cdxi6652m ^ cdxi6653m ^ cdxi6654m ^ cdxi6655m ^ cdxi6656m ^ cdxi6657m ^ cdxi6658m ^ cdxi6659m ^ cdxi6660m ^ cdxi6661m ^ cdxi6662m ^ cdxi6663m ^ cdxi6664m ^ cdxi6665m ^ cdxi6666m ^ cdxi6667m ^ cdxi6668m ^ cdxi6669m ^ cdxi6670m ^ cdxi6671m ^ cdxi6672m ^ cdxi6673m ^ cdxi6674m);
wire cdxi6676m = a1&cdxi6675m;
wire cdxi6677m = (reg_1_90);
wire cdxi6678m = (reg_1_100);
wire cdxi6679m = (reg_1_115);
wire cdxi6680m = reg_1_2&reg_1_5&reg_1_6&cdxi4738m;
wire cdxi6681m = reg_1_1&reg_1_5&reg_1_6&cdxi4795m;
wire cdxi6682m = reg_1_1&reg_1_2&cdxi5164m;
wire cdxi6683m = reg_1_1&reg_1_2&cdxi5165m;
wire cdxi6684m = reg_1_1&reg_1_2&cdxi5166m;
wire cdxi6685m = reg_1_5&cdxi5558m;
wire cdxi6686m = reg_1_2&reg_1_6&cdxi5004m;
wire cdxi6687m = reg_1_2&reg_1_5&reg_1_7&cdxi4905m;
wire cdxi6688m = reg_1_2&reg_1_5&reg_1_6&cdxi4737m;
wire cdxi6689m = reg_1_1&reg_1_6&cdxi5239m;
wire cdxi6690m = reg_1_1&reg_1_5&reg_1_7&cdxi4748m;
wire cdxi6691m = reg_1_1&reg_1_5&reg_1_6&cdxi4794m;
wire cdxi6692m = reg_1_1&reg_1_2&cdxi5167m;
wire cdxi6693m = reg_1_1&reg_1_2&cdxi5168m;
wire cdxi6694m = reg_1_1&reg_1_2&cdxi5169m;
wire cdxi6695m = reg_1_6&reg_1_7&cdxi5368m;
wire cdxi6696m = reg_1_5&cdxi5564m;
wire cdxi6697m = reg_1_5&cdxi5565m;
wire cdxi6698m = reg_1_2&reg_1_7&cdxi5515m;
wire cdxi6699m = reg_1_2&reg_1_6&cdxi5000m;
wire cdxi6700m = reg_1_2&reg_1_5&cdxi5551m;
wire cdxi6701m = reg_1_1&reg_1_7&cdxi5218m;
wire cdxi6702m = reg_1_1&reg_1_6&cdxi5235m;
wire cdxi6703m = reg_1_1&reg_1_5&cdxi5552m;
wire cdxi6704m = reg_1_1&reg_1_2&cdxi5163m;
wire cdxi6705m = reg_1_7&cdxi5516m;
wire cdxi6706m = reg_1_6&cdxi6470m;
wire cdxi6707m = reg_1_5&cdxi5553m;
wire cdxi6708m = reg_1_2&cdxi6677m;
wire cdxi6709m = reg_1_1&cdxi6678m;
wire cdxi6710m = (cdxi6680m ^ cdxi6681m ^ cdxi6682m ^ cdxi6683m ^ cdxi6684m ^ cdxi6685m ^ cdxi6686m ^ cdxi6687m ^ cdxi6688m ^ cdxi6689m ^ cdxi6690m ^ cdxi6691m ^ cdxi6692m ^ cdxi6693m ^ cdxi6694m ^ cdxi6695m ^ cdxi6696m ^ cdxi6697m ^ cdxi6698m ^ cdxi6699m ^ cdxi6700m ^ cdxi6701m ^ cdxi6702m ^ cdxi6703m ^ cdxi6704m ^ cdxi6705m ^ cdxi6706m ^ cdxi6707m ^ cdxi6708m ^ cdxi6709m ^ cdxi6679m);
wire cdxi6711m = reg_1_0&cdxi6710m;
wire cdxi6712m = cdxi4915m&cdxi5136m;
wire cdxi6713m = cdxi6712m&r0m;
wire cdxi6714m = cdxi5711m&cdxi4808m;
wire cdxi6715m = cdxi4874m&cdxi5137m;
wire cdxi6716m = cdxi4874m&cdxi5138m;
wire cdxi6717m = cdxi4874m&cdxi5139m;
wire cdxi6718m = cdxi5950m&r8m;
wire cdxi6719m = cdxi5083m&cdxi4977m;
wire cdxi6720m = cdxi5570m&r10m;
wire cdxi6721m = cdxi5779m&r11m;
wire cdxi6722m = cdxi4954m&cdxi5105m;
wire cdxi6723m = cdxi5463m&r19m;
wire cdxi6724m = cdxi5711m&r20m;
wire cdxi6725m = cdxi4874m&cdxi5140m;
wire cdxi6726m = cdxi4874m&cdxi5141m;
wire cdxi6727m = cdxi4874m&cdxi5142m;
wire cdxi6728m = cdxi5136m&r33m;
wire cdxi6729m = cdxi4973m&r34m;
wire cdxi6730m = cdxi4953m&r35m;
wire cdxi6731m = cdxi5101m&r37m;
wire cdxi6732m = cdxi5083m&r38m;
wire cdxi6733m = cdxi4915m&r40m;
wire cdxi6734m = cdxi4896m&r53m;
wire cdxi6735m = cdxi4954m&r54m;
wire cdxi6736m = cdxi4916m&r56m;
wire cdxi6737m = cdxi4874m&r59m;
wire cdxi6738m = cdxi4742m&r73m;
wire cdxi6739m = cdxi4762m&r74m;
wire cdxi6740m = cdxi4722m&r76m;
wire cdxi6741m = cdxi4711m&r79m;
wire cdxi6742m = cdxi4712m&r93m;
wire cdxi6743m = (cdxi108m ^ cdxi6713m ^ cdxi6714m ^ cdxi6715m ^ cdxi6716m ^ cdxi6717m ^ cdxi6718m ^ cdxi6719m ^ cdxi6720m ^ cdxi6721m ^ cdxi6722m ^ cdxi6723m ^ cdxi6724m ^ cdxi6725m ^ cdxi6726m ^ cdxi6727m ^ cdxi6728m ^ cdxi6729m ^ cdxi6730m ^ cdxi6731m ^ cdxi6732m ^ cdxi6733m ^ cdxi6734m ^ cdxi6735m ^ cdxi6736m ^ cdxi6737m ^ cdxi6738m ^ cdxi6739m ^ cdxi6740m ^ cdxi6741m ^ cdxi6742m);
wire cdxi6744m = a1&cdxi6743m;
wire cdxi6745m = (reg_1_116);
wire cdxi6746m = reg_1_3&reg_1_4&reg_1_5&reg_1_6&cdxi4664m;
wire cdxi6747m = reg_1_1&cdxi6169m;
wire cdxi6748m = reg_1_1&cdxi6170m;
wire cdxi6749m = reg_1_1&cdxi6171m;
wire cdxi6750m = reg_1_1&cdxi6172m;
wire cdxi6751m = reg_1_4&reg_1_5&reg_1_6&cdxi4717m;
wire cdxi6752m = reg_1_3&reg_1_5&cdxi4986m;
wire cdxi6753m = reg_1_3&reg_1_4&reg_1_6&cdxi4963m;
wire cdxi6754m = reg_1_3&reg_1_4&reg_1_5&cdxi4905m;
wire cdxi6755m = reg_1_1&cdxi6173m;
wire cdxi6756m = reg_1_1&cdxi6174m;
wire cdxi6757m = reg_1_1&cdxi6175m;
wire cdxi6758m = reg_1_1&cdxi6176m;
wire cdxi6759m = reg_1_1&cdxi6177m;
wire cdxi6760m = reg_1_1&cdxi6178m;
wire cdxi6761m = reg_1_5&cdxi5598m;
wire cdxi6762m = reg_1_4&reg_1_6&cdxi5369m;
wire cdxi6763m = reg_1_4&reg_1_5&cdxi5406m;
wire cdxi6764m = reg_1_3&reg_1_6&cdxi4964m;
wire cdxi6765m = reg_1_3&reg_1_5&cdxi4982m;
wire cdxi6766m = reg_1_3&reg_1_4&cdxi5515m;
wire cdxi6767m = reg_1_1&cdxi6179m;
wire cdxi6768m = reg_1_1&cdxi6180m;
wire cdxi6769m = reg_1_1&cdxi6181m;
wire cdxi6770m = reg_1_1&cdxi6182m;
wire cdxi6771m = reg_1_6&cdxi6262m;
wire cdxi6772m = reg_1_5&cdxi5587m;
wire cdxi6773m = reg_1_4&cdxi6400m;
wire cdxi6774m = reg_1_3&cdxi6538m;
wire cdxi6775m = reg_1_1&cdxi6168m;
wire cdxi6776m = (cdxi6746m ^ cdxi6747m ^ cdxi6748m ^ cdxi6749m ^ cdxi6750m ^ cdxi6751m ^ cdxi6752m ^ cdxi6753m ^ cdxi6754m ^ cdxi6755m ^ cdxi6756m ^ cdxi6757m ^ cdxi6758m ^ cdxi6759m ^ cdxi6760m ^ cdxi6761m ^ cdxi6762m ^ cdxi6763m ^ cdxi6764m ^ cdxi6765m ^ cdxi6766m ^ cdxi6767m ^ cdxi6768m ^ cdxi6769m ^ cdxi6770m ^ cdxi6771m ^ cdxi6772m ^ cdxi6773m ^ cdxi6774m ^ cdxi6775m ^ cdxi6745m);
wire cdxi6777m = reg_1_0&cdxi6776m;
wire cdxi6778m = cdxi4915m&cdxi4991m;
wire cdxi6779m = cdxi4916m&cdxi4991m;
wire cdxi6780m = cdxi4874m&cdxi5064m;
wire cdxi6781m = cdxi4915m&cdxi4992m;
wire cdxi6782m = cdxi4916m&cdxi5119m;
wire cdxi6783m = cdxi4874m&cdxi5292m;
wire cdxi6784m = cdxi4874m&cdxi5293m;
wire cdxi6785m = cdxi4874m&cdxi5294m;
wire cdxi6786m = cdxi4953m&cdxi4939m;
wire cdxi6787m = cdxi5640m&r9m;
wire cdxi6788m = cdxi4915m&cdxi4995m;
wire cdxi6789m = cdxi4915m&cdxi4996m;
wire cdxi6790m = cdxi4954m&cdxi5272m;
wire cdxi6791m = cdxi4916m&cdxi5122m;
wire cdxi6792m = cdxi4916m&cdxi5123m;
wire cdxi6793m = cdxi4874m&cdxi5295m;
wire cdxi6794m = cdxi4874m&cdxi5296m;
wire cdxi6795m = cdxi4874m&cdxi5297m;
wire cdxi6796m = cdxi4991m&r33m;
wire cdxi6797m = cdxi5064m&r34m;
wire cdxi6798m = cdxi4953m&r36m;
wire cdxi6799m = cdxi4934m&r37m;
wire cdxi6800m = cdxi5083m&r39m;
wire cdxi6801m = cdxi4915m&r41m;
wire cdxi6802m = cdxi4935m&r53m;
wire cdxi6803m = cdxi4954m&r55m;
wire cdxi6804m = cdxi4916m&r57m;
wire cdxi6805m = cdxi4874m&r60m;
wire cdxi6806m = cdxi4732m&r73m;
wire cdxi6807m = cdxi4762m&r75m;
wire cdxi6808m = cdxi4722m&r77m;
wire cdxi6809m = cdxi4711m&r80m;
wire cdxi6810m = cdxi4712m&r94m;
wire cdxi6811m = (cdxi109m ^ cdxi6781m ^ cdxi6782m ^ cdxi6783m ^ cdxi6784m ^ cdxi6785m ^ cdxi6786m ^ cdxi6787m ^ cdxi6788m ^ cdxi6789m ^ cdxi6790m ^ cdxi6791m ^ cdxi6792m ^ cdxi6793m ^ cdxi6794m ^ cdxi6795m ^ cdxi6796m ^ cdxi6797m ^ cdxi6798m ^ cdxi6799m ^ cdxi6800m ^ cdxi6801m ^ cdxi6802m ^ cdxi6803m ^ cdxi6804m ^ cdxi6805m ^ cdxi6806m ^ cdxi6807m ^ cdxi6808m ^ cdxi6809m ^ cdxi6810m);
wire cdxi6812m = a1&cdxi6811m;
wire cdxi6813m = (reg_1_117);
wire cdxi6814m = reg_1_3&cdxi5729m;
wire cdxi6815m = reg_1_1&cdxi6103m;
wire cdxi6816m = reg_1_1&cdxi6104m;
wire cdxi6817m = reg_1_1&cdxi6105m;
wire cdxi6818m = reg_1_1&cdxi6106m;
wire cdxi6819m = reg_1_4&cdxi5663m;
wire cdxi6820m = reg_1_3&cdxi5733m;
wire cdxi6821m = reg_1_3&cdxi5734m;
wire cdxi6822m = reg_1_3&cdxi5735m;
wire cdxi6823m = reg_1_1&cdxi6107m;
wire cdxi6824m = reg_1_1&cdxi6108m;
wire cdxi6825m = reg_1_1&cdxi6109m;
wire cdxi6826m = reg_1_1&cdxi6110m;
wire cdxi6827m = reg_1_1&cdxi6111m;
wire cdxi6828m = reg_1_1&cdxi6112m;
wire cdxi6829m = reg_1_5&cdxi5634m;
wire cdxi6830m = reg_1_4&cdxi5669m;
wire cdxi6831m = reg_1_4&cdxi5670m;
wire cdxi6832m = reg_1_3&cdxi5739m;
wire cdxi6833m = reg_1_3&cdxi5740m;
wire cdxi6834m = reg_1_3&cdxi5741m;
wire cdxi6835m = reg_1_1&cdxi6113m;
wire cdxi6836m = reg_1_1&cdxi6114m;
wire cdxi6837m = reg_1_1&cdxi6115m;
wire cdxi6838m = reg_1_1&cdxi6116m;
wire cdxi6839m = reg_1_7&cdxi6262m;
wire cdxi6840m = reg_1_5&cdxi5623m;
wire cdxi6841m = reg_1_4&cdxi5658m;
wire cdxi6842m = reg_1_3&cdxi5728m;
wire cdxi6843m = reg_1_1&cdxi6102m;
wire cdxi6844m = (cdxi6814m ^ cdxi6815m ^ cdxi6816m ^ cdxi6817m ^ cdxi6818m ^ cdxi6819m ^ cdxi6820m ^ cdxi6821m ^ cdxi6822m ^ cdxi6823m ^ cdxi6824m ^ cdxi6825m ^ cdxi6826m ^ cdxi6827m ^ cdxi6828m ^ cdxi6829m ^ cdxi6830m ^ cdxi6831m ^ cdxi6832m ^ cdxi6833m ^ cdxi6834m ^ cdxi6835m ^ cdxi6836m ^ cdxi6837m ^ cdxi6838m ^ cdxi6839m ^ cdxi6840m ^ cdxi6841m ^ cdxi6842m ^ cdxi6843m ^ cdxi6813m);
wire cdxi6845m = reg_1_0&cdxi6844m;
wire cdxi6846m = cdxi4953m&cdxi5154m;
wire cdxi6847m = cdxi5950m&cdxi4733m;
wire cdxi6848m = cdxi4954m&cdxi5250m;
wire cdxi6849m = cdxi4916m&cdxi5155m;
wire cdxi6850m = cdxi4916m&cdxi5156m;
wire cdxi6851m = cdxi4916m&cdxi5157m;
wire cdxi6852m = cdxi6017m&r9m;
wire cdxi6853m = cdxi4973m&cdxi4995m;
wire cdxi6854m = cdxi5710m&r11m;
wire cdxi6855m = cdxi5950m&r12m;
wire cdxi6856m = cdxi4896m&cdxi5295m;
wire cdxi6857m = cdxi4954m&cdxi5253m;
wire cdxi6858m = cdxi4954m&cdxi5254m;
wire cdxi6859m = cdxi4916m&cdxi5158m;
wire cdxi6860m = cdxi4916m&cdxi5159m;
wire cdxi6861m = cdxi4916m&cdxi5160m;
wire cdxi6862m = cdxi5154m&r37m;
wire cdxi6863m = cdxi4991m&r38m;
wire cdxi6864m = cdxi5136m&r39m;
wire cdxi6865m = cdxi5064m&r40m;
wire cdxi6866m = cdxi4973m&r41m;
wire cdxi6867m = cdxi4953m&r42m;
wire cdxi6868m = cdxi4935m&r59m;
wire cdxi6869m = cdxi4896m&r60m;
wire cdxi6870m = cdxi4954m&r61m;
wire cdxi6871m = cdxi4916m&r62m;
wire cdxi6872m = cdxi4732m&r79m;
wire cdxi6873m = cdxi4742m&r80m;
wire cdxi6874m = cdxi4762m&r81m;
wire cdxi6875m = cdxi4722m&r82m;
wire cdxi6876m = cdxi4712m&r97m;
wire cdxi6877m = (cdxi112m ^ cdxi6847m ^ cdxi6848m ^ cdxi6849m ^ cdxi6850m ^ cdxi6851m ^ cdxi6852m ^ cdxi6853m ^ cdxi6854m ^ cdxi6855m ^ cdxi6856m ^ cdxi6857m ^ cdxi6858m ^ cdxi6859m ^ cdxi6860m ^ cdxi6861m ^ cdxi6862m ^ cdxi6863m ^ cdxi6864m ^ cdxi6865m ^ cdxi6866m ^ cdxi6867m ^ cdxi6868m ^ cdxi6869m ^ cdxi6870m ^ cdxi6871m ^ cdxi6872m ^ cdxi6873m ^ cdxi6874m ^ cdxi6875m ^ cdxi6876m);
wire cdxi6878m = a1&cdxi6877m;
wire cdxi6879m = (reg_1_120);
wire cdxi6880m = reg_1_4&reg_1_5&reg_1_6&cdxi4738m;
wire cdxi6881m = reg_1_1&cdxi6208m;
wire cdxi6882m = reg_1_1&cdxi6209m;
wire cdxi6883m = reg_1_1&cdxi6210m;
wire cdxi6884m = reg_1_1&cdxi6211m;
wire cdxi6885m = reg_1_5&cdxi5767m;
wire cdxi6886m = reg_1_4&reg_1_6&cdxi5004m;
wire cdxi6887m = reg_1_4&reg_1_5&reg_1_7&cdxi4905m;
wire cdxi6888m = reg_1_4&reg_1_5&reg_1_6&cdxi4737m;
wire cdxi6889m = reg_1_1&cdxi6212m;
wire cdxi6890m = reg_1_1&cdxi6213m;
wire cdxi6891m = reg_1_1&cdxi6214m;
wire cdxi6892m = reg_1_1&cdxi6215m;
wire cdxi6893m = reg_1_1&cdxi6216m;
wire cdxi6894m = reg_1_1&cdxi6217m;
wire cdxi6895m = reg_1_6&cdxi5739m;
wire cdxi6896m = reg_1_5&cdxi5773m;
wire cdxi6897m = reg_1_5&cdxi5774m;
wire cdxi6898m = reg_1_4&reg_1_7&cdxi5515m;
wire cdxi6899m = reg_1_4&reg_1_6&cdxi5000m;
wire cdxi6900m = reg_1_4&reg_1_5&cdxi5551m;
wire cdxi6901m = reg_1_1&cdxi6218m;
wire cdxi6902m = reg_1_1&cdxi6219m;
wire cdxi6903m = reg_1_1&cdxi6220m;
wire cdxi6904m = reg_1_1&cdxi6221m;
wire cdxi6905m = reg_1_7&cdxi6538m;
wire cdxi6906m = reg_1_6&cdxi5728m;
wire cdxi6907m = reg_1_5&cdxi5762m;
wire cdxi6908m = reg_1_4&cdxi6677m;
wire cdxi6909m = reg_1_1&cdxi6207m;
wire cdxi6910m = (cdxi6880m ^ cdxi6881m ^ cdxi6882m ^ cdxi6883m ^ cdxi6884m ^ cdxi6885m ^ cdxi6886m ^ cdxi6887m ^ cdxi6888m ^ cdxi6889m ^ cdxi6890m ^ cdxi6891m ^ cdxi6892m ^ cdxi6893m ^ cdxi6894m ^ cdxi6895m ^ cdxi6896m ^ cdxi6897m ^ cdxi6898m ^ cdxi6899m ^ cdxi6900m ^ cdxi6901m ^ cdxi6902m ^ cdxi6903m ^ cdxi6904m ^ cdxi6905m ^ cdxi6906m ^ cdxi6907m ^ cdxi6908m ^ cdxi6909m ^ cdxi6879m);
wire cdxi6911m = reg_1_0&cdxi6910m;
wire cdxi6912m = cdxi4743m&cdxi5710m;
wire cdxi6913m = cdxi4873m&cdxi5064m;
wire cdxi6914m = cdxi4915m&cdxi5227m;
wire cdxi6915m = cdxi5780m&cdxi4753m;
wire cdxi6916m = cdxi4873m&cdxi5292m;
wire cdxi6917m = cdxi4873m&cdxi5293m;
wire cdxi6918m = cdxi4873m&cdxi5294m;
wire cdxi6919m = cdxi5710m&r13m;
wire cdxi6920m = cdxi5640m&r14m;
wire cdxi6921m = cdxi4915m&cdxi5230m;
wire cdxi6922m = cdxi4915m&cdxi5231m;
wire cdxi6923m = cdxi5883m&r18m;
wire cdxi6924m = cdxi5009m&cdxi5122m;
wire cdxi6925m = cdxi5780m&r21m;
wire cdxi6926m = cdxi4873m&cdxi5295m;
wire cdxi6927m = cdxi4873m&cdxi5296m;
wire cdxi6928m = cdxi4873m&cdxi5297m;
wire cdxi6929m = cdxi4991m&r43m;
wire cdxi6930m = cdxi5064m&r44m;
wire cdxi6931m = cdxi4953m&r46m;
wire cdxi6932m = cdxi4934m&r47m;
wire cdxi6933m = cdxi5083m&r49m;
wire cdxi6934m = cdxi4915m&r51m;
wire cdxi6935m = cdxi5065m&r53m;
wire cdxi6936m = cdxi5028m&r55m;
wire cdxi6937m = cdxi5009m&r57m;
wire cdxi6938m = cdxi4873m&r60m;
wire cdxi6939m = cdxi4732m&r83m;
wire cdxi6940m = cdxi4762m&r85m;
wire cdxi6941m = cdxi4722m&r87m;
wire cdxi6942m = cdxi4711m&r90m;
wire cdxi6943m = cdxi4743m&r94m;
wire cdxi6944m = (cdxi114m ^ cdxi6914m ^ cdxi6915m ^ cdxi6916m ^ cdxi6917m ^ cdxi6918m ^ cdxi6919m ^ cdxi6920m ^ cdxi6921m ^ cdxi6922m ^ cdxi6923m ^ cdxi6924m ^ cdxi6925m ^ cdxi6926m ^ cdxi6927m ^ cdxi6928m ^ cdxi6929m ^ cdxi6930m ^ cdxi6931m ^ cdxi6932m ^ cdxi6933m ^ cdxi6934m ^ cdxi6935m ^ cdxi6936m ^ cdxi6937m ^ cdxi6938m ^ cdxi6939m ^ cdxi6940m ^ cdxi6941m ^ cdxi6942m ^ cdxi6943m);
wire cdxi6945m = a1&cdxi6944m;
wire cdxi6946m = (reg_1_122);
wire cdxi6947m = reg_1_3&cdxi6001m;
wire cdxi6948m = reg_1_2&cdxi6103m;
wire cdxi6949m = reg_1_2&cdxi6104m;
wire cdxi6950m = reg_1_2&cdxi6105m;
wire cdxi6951m = reg_1_2&cdxi6106m;
wire cdxi6952m = reg_1_4&cdxi5905m;
wire cdxi6953m = reg_1_3&cdxi6005m;
wire cdxi6954m = reg_1_3&cdxi6006m;
wire cdxi6955m = reg_1_3&cdxi6007m;
wire cdxi6956m = reg_1_2&cdxi6107m;
wire cdxi6957m = reg_1_2&cdxi6108m;
wire cdxi6958m = reg_1_2&cdxi6109m;
wire cdxi6959m = reg_1_2&cdxi6110m;
wire cdxi6960m = reg_1_2&cdxi6111m;
wire cdxi6961m = reg_1_2&cdxi6112m;
wire cdxi6962m = reg_1_5&cdxi5842m;
wire cdxi6963m = reg_1_4&cdxi5911m;
wire cdxi6964m = reg_1_4&cdxi5912m;
wire cdxi6965m = reg_1_3&cdxi6011m;
wire cdxi6966m = reg_1_3&cdxi6012m;
wire cdxi6967m = reg_1_3&cdxi6013m;
wire cdxi6968m = reg_1_2&cdxi6113m;
wire cdxi6969m = reg_1_2&cdxi6114m;
wire cdxi6970m = reg_1_2&cdxi6115m;
wire cdxi6971m = reg_1_2&cdxi6116m;
wire cdxi6972m = reg_1_7&cdxi5797m;
wire cdxi6973m = reg_1_5&cdxi5831m;
wire cdxi6974m = reg_1_4&cdxi5900m;
wire cdxi6975m = reg_1_3&cdxi6000m;
wire cdxi6976m = reg_1_2&cdxi6102m;
wire cdxi6977m = (cdxi6947m ^ cdxi6948m ^ cdxi6949m ^ cdxi6950m ^ cdxi6951m ^ cdxi6952m ^ cdxi6953m ^ cdxi6954m ^ cdxi6955m ^ cdxi6956m ^ cdxi6957m ^ cdxi6958m ^ cdxi6959m ^ cdxi6960m ^ cdxi6961m ^ cdxi6962m ^ cdxi6963m ^ cdxi6964m ^ cdxi6965m ^ cdxi6966m ^ cdxi6967m ^ cdxi6968m ^ cdxi6969m ^ cdxi6970m ^ cdxi6971m ^ cdxi6972m ^ cdxi6973m ^ cdxi6974m ^ cdxi6975m ^ cdxi6976m ^ cdxi6946m);
wire cdxi6978m = reg_1_0&cdxi6977m;
wire cdxi6979m = cdxi4915m&cdxi5154m;
wire cdxi6980m = cdxi4873m&cdxi5154m;
wire cdxi6981m = cdxi5570m&cdxi4790m;
wire cdxi6982m = cdxi5462m&cdxi4753m;
wire cdxi6983m = cdxi4873m&cdxi5250m;
wire cdxi6984m = cdxi4873m&cdxi5251m;
wire cdxi6985m = cdxi4873m&cdxi5252m;
wire cdxi6986m = cdxi5745m&r13m;
wire cdxi6987m = cdxi5101m&cdxi5069m;
wire cdxi6988m = cdxi5604m&r16m;
wire cdxi6989m = cdxi5570m&r17m;
wire cdxi6990m = cdxi4895m&cdxi5272m;
wire cdxi6991m = cdxi5814m&r20m;
wire cdxi6992m = cdxi5462m&r21m;
wire cdxi6993m = cdxi4873m&cdxi5253m;
wire cdxi6994m = cdxi4873m&cdxi5254m;
wire cdxi6995m = cdxi4873m&cdxi5255m;
wire cdxi6996m = cdxi5154m&r43m;
wire cdxi6997m = cdxi5064m&r45m;
wire cdxi6998m = cdxi4973m&r46m;
wire cdxi6999m = cdxi4934m&r48m;
wire cdxi7000m = cdxi5101m&r49m;
wire cdxi7001m = cdxi4915m&r52m;
wire cdxi7002m = cdxi5065m&r54m;
wire cdxi7003m = cdxi4895m&r55m;
wire cdxi7004m = cdxi5009m&r58m;
wire cdxi7005m = cdxi4873m&r61m;
wire cdxi7006m = cdxi4732m&r84m;
wire cdxi7007m = cdxi4742m&r85m;
wire cdxi7008m = cdxi4722m&r88m;
wire cdxi7009m = cdxi4711m&r91m;
wire cdxi7010m = cdxi4743m&r95m;
wire cdxi7011m = (cdxi115m ^ cdxi6981m ^ cdxi6982m ^ cdxi6983m ^ cdxi6984m ^ cdxi6985m ^ cdxi6986m ^ cdxi6987m ^ cdxi6988m ^ cdxi6989m ^ cdxi6990m ^ cdxi6991m ^ cdxi6992m ^ cdxi6993m ^ cdxi6994m ^ cdxi6995m ^ cdxi6996m ^ cdxi6997m ^ cdxi6998m ^ cdxi6999m ^ cdxi7000m ^ cdxi7001m ^ cdxi7002m ^ cdxi7003m ^ cdxi7004m ^ cdxi7005m ^ cdxi7006m ^ cdxi7007m ^ cdxi7008m ^ cdxi7009m ^ cdxi7010m);
wire cdxi7012m = a1&cdxi7011m;
wire cdxi7013m = (reg_1_123);
wire cdxi7014m = reg_1_3&reg_1_4&reg_1_6&cdxi4795m;
wire cdxi7015m = reg_1_2&cdxi6136m;
wire cdxi7016m = reg_1_2&cdxi6137m;
wire cdxi7017m = reg_1_2&cdxi6138m;
wire cdxi7018m = reg_1_2&cdxi6139m;
wire cdxi7019m = reg_1_4&cdxi5938m;
wire cdxi7020m = reg_1_3&reg_1_6&cdxi5078m;
wire cdxi7021m = reg_1_3&reg_1_4&reg_1_7&cdxi4748m;
wire cdxi7022m = reg_1_3&reg_1_4&reg_1_6&cdxi4794m;
wire cdxi7023m = reg_1_2&cdxi6140m;
wire cdxi7024m = reg_1_2&cdxi6141m;
wire cdxi7025m = reg_1_2&cdxi6142m;
wire cdxi7026m = reg_1_2&cdxi6143m;
wire cdxi7027m = reg_1_2&cdxi6144m;
wire cdxi7028m = reg_1_2&cdxi6145m;
wire cdxi7029m = reg_1_6&cdxi5842m;
wire cdxi7030m = reg_1_4&cdxi5944m;
wire cdxi7031m = reg_1_4&cdxi5945m;
wire cdxi7032m = reg_1_3&reg_1_7&cdxi5055m;
wire cdxi7033m = reg_1_3&reg_1_6&cdxi5074m;
wire cdxi7034m = reg_1_3&reg_1_4&cdxi5552m;
wire cdxi7035m = reg_1_2&cdxi6146m;
wire cdxi7036m = reg_1_2&cdxi6147m;
wire cdxi7037m = reg_1_2&cdxi6148m;
wire cdxi7038m = reg_1_2&cdxi6149m;
wire cdxi7039m = reg_1_7&cdxi6067m;
wire cdxi7040m = reg_1_6&cdxi5831m;
wire cdxi7041m = reg_1_4&cdxi5933m;
wire cdxi7042m = reg_1_3&cdxi6609m;
wire cdxi7043m = reg_1_2&cdxi6135m;
wire cdxi7044m = (cdxi7014m ^ cdxi7015m ^ cdxi7016m ^ cdxi7017m ^ cdxi7018m ^ cdxi7019m ^ cdxi7020m ^ cdxi7021m ^ cdxi7022m ^ cdxi7023m ^ cdxi7024m ^ cdxi7025m ^ cdxi7026m ^ cdxi7027m ^ cdxi7028m ^ cdxi7029m ^ cdxi7030m ^ cdxi7031m ^ cdxi7032m ^ cdxi7033m ^ cdxi7034m ^ cdxi7035m ^ cdxi7036m ^ cdxi7037m ^ cdxi7038m ^ cdxi7039m ^ cdxi7040m ^ cdxi7041m ^ cdxi7042m ^ cdxi7043m ^ cdxi7013m);
wire cdxi7045m = reg_1_0&cdxi7044m;
wire cdxi7046m = cdxi5950m&cdxi4790m;
wire cdxi7047m = cdxi5028m&cdxi5250m;
wire cdxi7048m = cdxi5462m&cdxi4781m;
wire cdxi7049m = cdxi5780m&cdxi4850m;
wire cdxi7050m = cdxi5780m&cdxi4851m;
wire cdxi7051m = cdxi5136m&cdxi5069m;
wire cdxi7052m = cdxi4973m&cdxi5230m;
wire cdxi7053m = cdxi5710m&r16m;
wire cdxi7054m = cdxi5950m&r17m;
wire cdxi7055m = cdxi4895m&cdxi5295m;
wire cdxi7056m = cdxi5883m&r23m;
wire cdxi7057m = cdxi5028m&cdxi5254m;
wire cdxi7058m = cdxi5009m&cdxi5158m;
wire cdxi7059m = cdxi5462m&r26m;
wire cdxi7060m = cdxi5780m&r27m;
wire cdxi7061m = cdxi5154m&r47m;
wire cdxi7062m = cdxi4991m&r48m;
wire cdxi7063m = cdxi5136m&r49m;
wire cdxi7064m = cdxi5064m&r50m;
wire cdxi7065m = cdxi4973m&r51m;
wire cdxi7066m = cdxi4953m&r52m;
wire cdxi7067m = cdxi5065m&r59m;
wire cdxi7068m = cdxi4895m&r60m;
wire cdxi7069m = cdxi5028m&r61m;
wire cdxi7070m = cdxi5009m&r62m;
wire cdxi7071m = cdxi4732m&r89m;
wire cdxi7072m = cdxi4742m&r90m;
wire cdxi7073m = cdxi4762m&r91m;
wire cdxi7074m = cdxi4722m&r92m;
wire cdxi7075m = cdxi4743m&r97m;
wire cdxi7076m = (cdxi117m ^ cdxi7046m ^ cdxi7047m ^ cdxi7048m ^ cdxi7049m ^ cdxi7050m ^ cdxi7051m ^ cdxi7052m ^ cdxi7053m ^ cdxi7054m ^ cdxi7055m ^ cdxi7056m ^ cdxi7057m ^ cdxi7058m ^ cdxi7059m ^ cdxi7060m ^ cdxi7061m ^ cdxi7062m ^ cdxi7063m ^ cdxi7064m ^ cdxi7065m ^ cdxi7066m ^ cdxi7067m ^ cdxi7068m ^ cdxi7069m ^ cdxi7070m ^ cdxi7071m ^ cdxi7072m ^ cdxi7073m ^ cdxi7074m ^ cdxi7075m);
wire cdxi7077m = a1&cdxi7076m;
wire cdxi7078m = (reg_1_125);
wire cdxi7079m = reg_1_4&reg_1_5&reg_1_6&cdxi4795m;
wire cdxi7080m = reg_1_2&cdxi6208m;
wire cdxi7081m = reg_1_2&cdxi6209m;
wire cdxi7082m = reg_1_2&cdxi6210m;
wire cdxi7083m = reg_1_2&cdxi6211m;
wire cdxi7084m = reg_1_5&reg_1_6&cdxi5078m;
wire cdxi7085m = reg_1_4&reg_1_6&cdxi5239m;
wire cdxi7086m = reg_1_4&reg_1_5&reg_1_7&cdxi4748m;
wire cdxi7087m = reg_1_4&reg_1_5&reg_1_6&cdxi4794m;
wire cdxi7088m = reg_1_2&cdxi6212m;
wire cdxi7089m = reg_1_2&cdxi6213m;
wire cdxi7090m = reg_1_2&cdxi6214m;
wire cdxi7091m = reg_1_2&cdxi6215m;
wire cdxi7092m = reg_1_2&cdxi6216m;
wire cdxi7093m = reg_1_2&cdxi6217m;
wire cdxi7094m = reg_1_6&cdxi6011m;
wire cdxi7095m = reg_1_5&reg_1_7&cdxi5055m;
wire cdxi7096m = reg_1_5&reg_1_6&cdxi5074m;
wire cdxi7097m = reg_1_4&reg_1_7&cdxi5218m;
wire cdxi7098m = reg_1_4&reg_1_6&cdxi5235m;
wire cdxi7099m = reg_1_4&reg_1_5&cdxi5552m;
wire cdxi7100m = reg_1_2&cdxi6218m;
wire cdxi7101m = reg_1_2&cdxi6219m;
wire cdxi7102m = reg_1_2&cdxi6220m;
wire cdxi7103m = reg_1_2&cdxi6221m;
wire cdxi7104m = reg_1_7&cdxi5967m;
wire cdxi7105m = reg_1_6&cdxi6000m;
wire cdxi7106m = reg_1_5&cdxi6609m;
wire cdxi7107m = reg_1_4&cdxi6678m;
wire cdxi7108m = reg_1_2&cdxi6207m;
wire cdxi7109m = (cdxi7079m ^ cdxi7080m ^ cdxi7081m ^ cdxi7082m ^ cdxi7083m ^ cdxi7084m ^ cdxi7085m ^ cdxi7086m ^ cdxi7087m ^ cdxi7088m ^ cdxi7089m ^ cdxi7090m ^ cdxi7091m ^ cdxi7092m ^ cdxi7093m ^ cdxi7094m ^ cdxi7095m ^ cdxi7096m ^ cdxi7097m ^ cdxi7098m ^ cdxi7099m ^ cdxi7100m ^ cdxi7101m ^ cdxi7102m ^ cdxi7103m ^ cdxi7104m ^ cdxi7105m ^ cdxi7106m ^ cdxi7107m ^ cdxi7108m ^ cdxi7078m);
wire cdxi7110m = reg_1_0&cdxi7109m;
wire cdxi7111m = cdxi5083m&cdxi5154m;
wire cdxi7112m = cdxi5950m&cdxi4753m;
wire cdxi7113m = cdxi5083m&cdxi5250m;
wire cdxi7114m = cdxi4915m&cdxi5155m;
wire cdxi7115m = cdxi4915m&cdxi5156m;
wire cdxi7116m = cdxi4915m&cdxi5157m;
wire cdxi7117m = cdxi5136m&cdxi5272m;
wire cdxi7118m = cdxi4973m&cdxi5122m;
wire cdxi7119m = cdxi5710m&r20m;
wire cdxi7120m = cdxi5950m&r21m;
wire cdxi7121m = cdxi5101m&cdxi5295m;
wire cdxi7122m = cdxi5640m&r23m;
wire cdxi7123m = cdxi5083m&cdxi5254m;
wire cdxi7124m = cdxi4915m&cdxi5158m;
wire cdxi7125m = cdxi4915m&cdxi5159m;
wire cdxi7126m = cdxi4915m&cdxi5160m;
wire cdxi7127m = cdxi5154m&r53m;
wire cdxi7128m = cdxi4991m&r54m;
wire cdxi7129m = cdxi5136m&r55m;
wire cdxi7130m = cdxi5064m&r56m;
wire cdxi7131m = cdxi4973m&r57m;
wire cdxi7132m = cdxi4953m&r58m;
wire cdxi7133m = cdxi4934m&r59m;
wire cdxi7134m = cdxi5101m&r60m;
wire cdxi7135m = cdxi5083m&r61m;
wire cdxi7136m = cdxi4915m&r62m;
wire cdxi7137m = cdxi4732m&r93m;
wire cdxi7138m = cdxi4742m&r94m;
wire cdxi7139m = cdxi4762m&r95m;
wire cdxi7140m = cdxi4722m&r96m;
wire cdxi7141m = cdxi4711m&r97m;
wire cdxi7142m = (cdxi118m ^ cdxi7112m ^ cdxi7113m ^ cdxi7114m ^ cdxi7115m ^ cdxi7116m ^ cdxi7117m ^ cdxi7118m ^ cdxi7119m ^ cdxi7120m ^ cdxi7121m ^ cdxi7122m ^ cdxi7123m ^ cdxi7124m ^ cdxi7125m ^ cdxi7126m ^ cdxi7127m ^ cdxi7128m ^ cdxi7129m ^ cdxi7130m ^ cdxi7131m ^ cdxi7132m ^ cdxi7133m ^ cdxi7134m ^ cdxi7135m ^ cdxi7136m ^ cdxi7137m ^ cdxi7138m ^ cdxi7139m ^ cdxi7140m ^ cdxi7141m);
wire cdxi7143m = a1&cdxi7142m;
wire cdxi7144m = (reg_1_126);
wire cdxi7145m = reg_1_4&cdxi6035m;
wire cdxi7146m = reg_1_3&cdxi6208m;
wire cdxi7147m = reg_1_3&cdxi6209m;
wire cdxi7148m = reg_1_3&cdxi6210m;
wire cdxi7149m = reg_1_3&cdxi6211m;
wire cdxi7150m = reg_1_5&cdxi6140m;
wire cdxi7151m = reg_1_4&cdxi6039m;
wire cdxi7152m = reg_1_4&cdxi6040m;
wire cdxi7153m = reg_1_4&cdxi6041m;
wire cdxi7154m = reg_1_3&cdxi6212m;
wire cdxi7155m = reg_1_3&cdxi6213m;
wire cdxi7156m = reg_1_3&cdxi6214m;
wire cdxi7157m = reg_1_3&cdxi6215m;
wire cdxi7158m = reg_1_3&cdxi6216m;
wire cdxi7159m = reg_1_3&cdxi6217m;
wire cdxi7160m = reg_1_6&cdxi6113m;
wire cdxi7161m = reg_1_5&cdxi6146m;
wire cdxi7162m = reg_1_5&cdxi6147m;
wire cdxi7163m = reg_1_4&cdxi6045m;
wire cdxi7164m = reg_1_4&cdxi6046m;
wire cdxi7165m = reg_1_4&cdxi6047m;
wire cdxi7166m = reg_1_3&cdxi6218m;
wire cdxi7167m = reg_1_3&cdxi6219m;
wire cdxi7168m = reg_1_3&cdxi6220m;
wire cdxi7169m = reg_1_3&cdxi6221m;
wire cdxi7170m = reg_1_7&cdxi6168m;
wire cdxi7171m = reg_1_6&cdxi6102m;
wire cdxi7172m = reg_1_5&cdxi6135m;
wire cdxi7173m = reg_1_4&cdxi6034m;
wire cdxi7174m = reg_1_3&cdxi6207m;
wire cdxi7175m = (cdxi7145m ^ cdxi7146m ^ cdxi7147m ^ cdxi7148m ^ cdxi7149m ^ cdxi7150m ^ cdxi7151m ^ cdxi7152m ^ cdxi7153m ^ cdxi7154m ^ cdxi7155m ^ cdxi7156m ^ cdxi7157m ^ cdxi7158m ^ cdxi7159m ^ cdxi7160m ^ cdxi7161m ^ cdxi7162m ^ cdxi7163m ^ cdxi7164m ^ cdxi7165m ^ cdxi7166m ^ cdxi7167m ^ cdxi7168m ^ cdxi7169m ^ cdxi7170m ^ cdxi7171m ^ cdxi7172m ^ cdxi7173m ^ cdxi7174m ^ cdxi7144m);
wire cdxi7176m = reg_1_0&cdxi7175m;
wire cdxi7177m = cdxi4712m&cdxi6944m;
wire cdxi7178m = reg_1_1&cdxi6977m;
wire cdxi7179m = cdxi4712m&cdxi7011m;
wire cdxi7180m = reg_1_1&cdxi7044m;
wire cdxi7181m = cdxi5848m&cdxi4790m;
wire cdxi7182m = cdxi5497m&cdxi4753m;
wire cdxi7183m = cdxi4873m&cdxi5155m;
wire cdxi7184m = cdxi4873m&cdxi5156m;
wire cdxi7185m = cdxi4873m&cdxi5157m;
wire cdxi7186m = cdxi6017m&r13m;
wire cdxi7187m = cdxi5101m&cdxi5230m;
wire cdxi7188m = cdxi5640m&r16m;
wire cdxi7189m = cdxi5848m&r17m;
wire cdxi7190m = cdxi4895m&cdxi5122m;
wire cdxi7191m = cdxi5883m&r20m;
wire cdxi7192m = cdxi5497m&r21m;
wire cdxi7193m = cdxi4873m&cdxi5158m;
wire cdxi7194m = cdxi4873m&cdxi5159m;
wire cdxi7195m = cdxi4873m&cdxi5160m;
wire cdxi7196m = cdxi5154m&r44m;
wire cdxi7197m = cdxi4991m&r45m;
wire cdxi7198m = cdxi5136m&r46m;
wire cdxi7199m = cdxi4934m&r50m;
wire cdxi7200m = cdxi5101m&r51m;
wire cdxi7201m = cdxi5083m&r52m;
wire cdxi7202m = cdxi5065m&r56m;
wire cdxi7203m = cdxi4895m&r57m;
wire cdxi7204m = cdxi5028m&r58m;
wire cdxi7205m = cdxi4873m&r62m;
wire cdxi7206m = cdxi4732m&r86m;
wire cdxi7207m = cdxi4742m&r87m;
wire cdxi7208m = cdxi4762m&r88m;
wire cdxi7209m = cdxi4711m&r92m;
wire cdxi7210m = cdxi4743m&r96m;
wire cdxi7211m = (cdxi116m ^ cdxi7181m ^ cdxi7182m ^ cdxi7183m ^ cdxi7184m ^ cdxi7185m ^ cdxi7186m ^ cdxi7187m ^ cdxi7188m ^ cdxi7189m ^ cdxi7190m ^ cdxi7191m ^ cdxi7192m ^ cdxi7193m ^ cdxi7194m ^ cdxi7195m ^ cdxi7196m ^ cdxi7197m ^ cdxi7198m ^ cdxi7199m ^ cdxi7200m ^ cdxi7201m ^ cdxi7202m ^ cdxi7203m ^ cdxi7204m ^ cdxi7205m ^ cdxi7206m ^ cdxi7207m ^ cdxi7208m ^ cdxi7209m ^ cdxi7210m);
wire cdxi7212m = cdxi4712m&cdxi7211m;
wire cdxi7213m = (reg_1_124);
wire cdxi7214m = reg_1_3&reg_1_5&reg_1_6&cdxi4795m;
wire cdxi7215m = reg_1_2&cdxi6035m;
wire cdxi7216m = reg_1_2&cdxi6036m;
wire cdxi7217m = reg_1_2&cdxi6037m;
wire cdxi7218m = reg_1_2&cdxi6038m;
wire cdxi7219m = reg_1_5&cdxi5938m;
wire cdxi7220m = reg_1_3&reg_1_6&cdxi5239m;
wire cdxi7221m = reg_1_3&reg_1_5&reg_1_7&cdxi4748m;
wire cdxi7222m = reg_1_3&reg_1_5&reg_1_6&cdxi4794m;
wire cdxi7223m = reg_1_2&cdxi6039m;
wire cdxi7224m = reg_1_2&cdxi6040m;
wire cdxi7225m = reg_1_2&cdxi6041m;
wire cdxi7226m = reg_1_2&cdxi6042m;
wire cdxi7227m = reg_1_2&cdxi6043m;
wire cdxi7228m = reg_1_2&cdxi6044m;
wire cdxi7229m = reg_1_6&cdxi5911m;
wire cdxi7230m = reg_1_5&cdxi5944m;
wire cdxi7231m = reg_1_5&cdxi5945m;
wire cdxi7232m = reg_1_3&reg_1_7&cdxi5218m;
wire cdxi7233m = reg_1_3&reg_1_6&cdxi5235m;
wire cdxi7234m = reg_1_3&reg_1_5&cdxi5552m;
wire cdxi7235m = reg_1_2&cdxi6045m;
wire cdxi7236m = reg_1_2&cdxi6046m;
wire cdxi7237m = reg_1_2&cdxi6047m;
wire cdxi7238m = reg_1_2&cdxi6048m;
wire cdxi7239m = reg_1_7&cdxi5866m;
wire cdxi7240m = reg_1_6&cdxi5900m;
wire cdxi7241m = reg_1_5&cdxi5933m;
wire cdxi7242m = reg_1_3&cdxi6678m;
wire cdxi7243m = reg_1_2&cdxi6034m;
wire cdxi7244m = (cdxi7214m ^ cdxi7215m ^ cdxi7216m ^ cdxi7217m ^ cdxi7218m ^ cdxi7219m ^ cdxi7220m ^ cdxi7221m ^ cdxi7222m ^ cdxi7223m ^ cdxi7224m ^ cdxi7225m ^ cdxi7226m ^ cdxi7227m ^ cdxi7228m ^ cdxi7229m ^ cdxi7230m ^ cdxi7231m ^ cdxi7232m ^ cdxi7233m ^ cdxi7234m ^ cdxi7235m ^ cdxi7236m ^ cdxi7237m ^ cdxi7238m ^ cdxi7239m ^ cdxi7240m ^ cdxi7241m ^ cdxi7242m ^ cdxi7243m ^ cdxi7213m);
wire cdxi7245m = reg_1_1&cdxi7244m;
wire cdxi7246m = cdxi4712m&cdxi7142m;
wire cdxi7247m = reg_1_1&cdxi7175m;
wire cdxi7248m = cdxi4873m&cdxi5745m;
wire cdxi7249m = cdxi4874m&cdxi5745m;
wire cdxi7250m = cdxi4875m&cdxi5745m;
wire cdxi7251m = cdxi5314m&cdxi5154m;
wire cdxi7252m = cdxi5314m&cdxi5064m;
wire cdxi7253m = cdxi5314m&cdxi4973m;
wire cdxi7254m = cdxi4874m&cdxi5154m;
wire cdxi7255m = cdxi4873m&cdxi5746m;
wire cdxi7256m = cdxi6297m&cdxi4790m;
wire cdxi7257m = cdxi4875m&cdxi6119m;
wire cdxi7258m = cdxi5314m&cdxi5250m;
wire cdxi7259m = cdxi5314m&cdxi5251m;
wire cdxi7260m = cdxi5314m&cdxi5252m;
wire cdxi7261m = cdxi4915m&cdxi5539m;
wire cdxi7262m = cdxi5462m&cdxi4939m;
wire cdxi7263m = cdxi4873m&cdxi5750m;
wire cdxi7264m = cdxi4873m&cdxi5751m;
wire cdxi7265m = cdxi4873m&cdxi5752m;
wire cdxi7266m = cdxi4916m&cdxi5921m;
wire cdxi7267m = cdxi5388m&cdxi5069m;
wire cdxi7268m = cdxi6780m&r16m;
wire cdxi7269m = cdxi6297m&r17m;
wire cdxi7270m = cdxi4875m&cdxi6123m;
wire cdxi7271m = cdxi4875m&cdxi6124m;
wire cdxi7272m = cdxi4875m&cdxi6125m;
wire cdxi7273m = cdxi5314m&cdxi5253m;
wire cdxi7274m = cdxi5314m&cdxi5254m;
wire cdxi7275m = cdxi5314m&cdxi5255m;
wire cdxi7276m = cdxi4973m&cdxi5437m;
wire cdxi7277m = cdxi5675m&r29m;
wire cdxi7278m = cdxi4915m&cdxi5545m;
wire cdxi7279m = cdxi4915m&cdxi5546m;
wire cdxi7280m = cdxi5533m&r33m;
wire cdxi7281m = cdxi5009m&cdxi5686m;
wire cdxi7282m = cdxi5462m&r36m;
wire cdxi7283m = cdxi5424m&r38m;
wire cdxi7284m = cdxi5387m&r39m;
wire cdxi7285m = cdxi5311m&r42m;
wire cdxi7286m = cdxi5534m&r43m;
wire cdxi7287m = cdxi5605m&r45m;
wire cdxi7288m = cdxi5463m&r46m;
wire cdxi7289m = cdxi5425m&r48m;
wire cdxi7290m = cdxi5388m&r49m;
wire cdxi7291m = cdxi5312m&r52m;
wire cdxi7292m = cdxi5426m&r54m;
wire cdxi7293m = cdxi5389m&r55m;
wire cdxi7294m = cdxi5313m&r58m;
wire cdxi7295m = cdxi5314m&r61m;
wire cdxi7296m = cdxi5154m&r63m;
wire cdxi7297m = cdxi5064m&r65m;
wire cdxi7298m = cdxi4973m&r66m;
wire cdxi7299m = cdxi4934m&r68m;
wire cdxi7300m = cdxi5101m&r69m;
wire cdxi7301m = cdxi4915m&r72m;
wire cdxi7302m = cdxi5065m&r74m;
wire cdxi7303m = cdxi4895m&r75m;
wire cdxi7304m = cdxi5009m&r78m;
wire cdxi7305m = cdxi4873m&r81m;
wire cdxi7306m = cdxi4935m&r84m;
wire cdxi7307m = cdxi4896m&r85m;
wire cdxi7308m = cdxi4916m&r88m;
wire cdxi7309m = cdxi4874m&r91m;
wire cdxi7310m = cdxi4875m&r95m;
wire cdxi7311m = cdxi4732m&r99m;
wire cdxi7312m = cdxi4742m&r100m;
wire cdxi7313m = cdxi4722m&r103m;
wire cdxi7314m = cdxi4711m&r106m;
wire cdxi7315m = cdxi4743m&r110m;
wire cdxi7316m = cdxi4712m&r115m;
wire cdxi7317m = (cdxi121m ^ cdxi7255m ^ cdxi7256m ^ cdxi7257m ^ cdxi7258m ^ cdxi7259m ^ cdxi7260m ^ cdxi7261m ^ cdxi7262m ^ cdxi7263m ^ cdxi7264m ^ cdxi7265m ^ cdxi7266m ^ cdxi7267m ^ cdxi7268m ^ cdxi7269m ^ cdxi7270m ^ cdxi7271m ^ cdxi7272m ^ cdxi7273m ^ cdxi7274m ^ cdxi7275m ^ cdxi7276m ^ cdxi7277m ^ cdxi7278m ^ cdxi7279m ^ cdxi7280m ^ cdxi7281m ^ cdxi7282m ^ cdxi7283m ^ cdxi7284m ^ cdxi7285m ^ cdxi7286m ^ cdxi7287m ^ cdxi7288m ^ cdxi7289m ^ cdxi7290m ^ cdxi7291m ^ cdxi7292m ^ cdxi7293m ^ cdxi7294m ^ cdxi7295m ^ cdxi7296m ^ cdxi7297m ^ cdxi7298m ^ cdxi7299m ^ cdxi7300m ^ cdxi7301m ^ cdxi7302m ^ cdxi7303m ^ cdxi7304m ^ cdxi7305m ^ cdxi7306m ^ cdxi7307m ^ cdxi7308m ^ cdxi7309m ^ cdxi7310m ^ cdxi7311m ^ cdxi7312m ^ cdxi7313m ^ cdxi7314m ^ cdxi7315m ^ cdxi7316m);
wire cdxi7318m = a1&cdxi7317m;
wire cdxi7319m = (reg_1_108);
wire cdxi7320m = (reg_1_111);
wire cdxi7321m = (reg_1_118);
wire cdxi7322m = (reg_1_129);
wire cdxi7323m = reg_1_2&reg_1_3&cdxi5763m;
wire cdxi7324m = reg_1_1&cdxi7014m;
wire cdxi7325m = reg_1_1&cdxi7015m;
wire cdxi7326m = reg_1_1&cdxi7016m;
wire cdxi7327m = reg_1_1&cdxi7017m;
wire cdxi7328m = reg_1_1&cdxi7018m;
wire cdxi7329m = reg_1_3&cdxi6616m;
wire cdxi7330m = reg_1_2&reg_1_4&cdxi5698m;
wire cdxi7331m = reg_1_2&reg_1_3&cdxi5767m;
wire cdxi7332m = reg_1_2&reg_1_3&cdxi5768m;
wire cdxi7333m = reg_1_2&reg_1_3&cdxi5769m;
wire cdxi7334m = reg_1_1&cdxi7019m;
wire cdxi7335m = reg_1_1&cdxi7020m;
wire cdxi7336m = reg_1_1&cdxi7021m;
wire cdxi7337m = reg_1_1&cdxi7022m;
wire cdxi7338m = reg_1_1&cdxi7023m;
wire cdxi7339m = reg_1_1&cdxi7024m;
wire cdxi7340m = reg_1_1&cdxi7025m;
wire cdxi7341m = reg_1_1&cdxi7026m;
wire cdxi7342m = reg_1_1&cdxi7027m;
wire cdxi7343m = reg_1_1&cdxi7028m;
wire cdxi7344m = reg_1_4&reg_1_6&cdxi5456m;
wire cdxi7345m = reg_1_3&cdxi6626m;
wire cdxi7346m = reg_1_3&cdxi6627m;
wire cdxi7347m = reg_1_3&cdxi6628m;
wire cdxi7348m = reg_1_2&reg_1_6&cdxi5634m;
wire cdxi7349m = reg_1_2&reg_1_4&cdxi5704m;
wire cdxi7350m = reg_1_2&reg_1_4&cdxi5705m;
wire cdxi7351m = reg_1_2&reg_1_3&cdxi5773m;
wire cdxi7352m = reg_1_2&reg_1_3&cdxi5774m;
wire cdxi7353m = reg_1_2&reg_1_3&cdxi5775m;
wire cdxi7354m = reg_1_1&cdxi7029m;
wire cdxi7355m = reg_1_1&cdxi7030m;
wire cdxi7356m = reg_1_1&cdxi7031m;
wire cdxi7357m = reg_1_1&cdxi7032m;
wire cdxi7358m = reg_1_1&cdxi7033m;
wire cdxi7359m = reg_1_1&cdxi7034m;
wire cdxi7360m = reg_1_1&cdxi7035m;
wire cdxi7361m = reg_1_1&cdxi7036m;
wire cdxi7362m = reg_1_1&cdxi7037m;
wire cdxi7363m = reg_1_1&cdxi7038m;
wire cdxi7364m = reg_1_6&reg_1_7&cdxi5332m;
wire cdxi7365m = reg_1_4&reg_1_7&cdxi5407m;
wire cdxi7366m = reg_1_4&reg_1_6&cdxi5445m;
wire cdxi7367m = reg_1_3&cdxi6636m;
wire cdxi7368m = reg_1_3&cdxi6637m;
wire cdxi7369m = reg_1_3&cdxi6638m;
wire cdxi7370m = reg_1_2&reg_1_7&cdxi5587m;
wire cdxi7371m = reg_1_2&reg_1_6&cdxi5623m;
wire cdxi7372m = reg_1_2&reg_1_4&cdxi5693m;
wire cdxi7373m = reg_1_2&reg_1_3&cdxi5762m;
wire cdxi7374m = reg_1_1&cdxi7039m;
wire cdxi7375m = reg_1_1&cdxi7040m;
wire cdxi7376m = reg_1_1&cdxi7041m;
wire cdxi7377m = reg_1_1&cdxi7042m;
wire cdxi7378m = reg_1_1&cdxi7043m;
wire cdxi7379m = reg_1_7&cdxi6332m;
wire cdxi7380m = reg_1_6&cdxi7319m;
wire cdxi7381m = reg_1_4&cdxi7320m;
wire cdxi7382m = reg_1_3&cdxi6610m;
wire cdxi7383m = reg_1_2&cdxi7321m;
wire cdxi7384m = reg_1_1&cdxi7013m;
wire cdxi7385m = (cdxi7323m ^ cdxi7324m ^ cdxi7325m ^ cdxi7326m ^ cdxi7327m ^ cdxi7328m ^ cdxi7329m ^ cdxi7330m ^ cdxi7331m ^ cdxi7332m ^ cdxi7333m ^ cdxi7334m ^ cdxi7335m ^ cdxi7336m ^ cdxi7337m ^ cdxi7338m ^ cdxi7339m ^ cdxi7340m ^ cdxi7341m ^ cdxi7342m ^ cdxi7343m ^ cdxi7344m ^ cdxi7345m ^ cdxi7346m ^ cdxi7347m ^ cdxi7348m ^ cdxi7349m ^ cdxi7350m ^ cdxi7351m ^ cdxi7352m ^ cdxi7353m ^ cdxi7354m ^ cdxi7355m ^ cdxi7356m ^ cdxi7357m ^ cdxi7358m ^ cdxi7359m ^ cdxi7360m ^ cdxi7361m ^ cdxi7362m ^ cdxi7363m ^ cdxi7364m ^ cdxi7365m ^ cdxi7366m ^ cdxi7367m ^ cdxi7368m ^ cdxi7369m ^ cdxi7370m ^ cdxi7371m ^ cdxi7372m ^ cdxi7373m ^ cdxi7374m ^ cdxi7375m ^ cdxi7376m ^ cdxi7377m ^ cdxi7378m ^ cdxi7379m ^ cdxi7380m ^ cdxi7381m ^ cdxi7382m ^ cdxi7383m ^ cdxi7384m ^ cdxi7322m);
wire cdxi7386m = reg_1_0&cdxi7385m;
wire cdxi7387m = cdxi4873m&cdxi6017m;
wire cdxi7388m = cdxi4874m&cdxi6017m;
wire cdxi7389m = cdxi4875m&cdxi6017m;
wire cdxi7390m = cdxi5314m&cdxi4991m;
wire cdxi7391m = cdxi5314m&cdxi5136m;
wire cdxi7392m = cdxi6365m&cdxi4733m;
wire cdxi7393m = cdxi6366m&cdxi4790m;
wire cdxi7394m = cdxi4875m&cdxi6018m;
wire cdxi7395m = cdxi5314m&cdxi5155m;
wire cdxi7396m = cdxi5314m&cdxi5156m;
wire cdxi7397m = cdxi5314m&cdxi5157m;
wire cdxi7398m = cdxi5083m&cdxi5539m;
wire cdxi7399m = cdxi5497m&cdxi4939m;
wire cdxi7400m = cdxi5387m&cdxi4995m;
wire cdxi7401m = cdxi6434m&r11m;
wire cdxi7402m = cdxi6365m&r12m;
wire cdxi7403m = cdxi4954m&cdxi5921m;
wire cdxi7404m = cdxi7254m&r15m;
wire cdxi7405m = cdxi6435m&r16m;
wire cdxi7406m = cdxi6366m&r17m;
wire cdxi7407m = cdxi5389m&cdxi5122m;
wire cdxi7408m = cdxi4875m&cdxi6023m;
wire cdxi7409m = cdxi4875m&cdxi6024m;
wire cdxi7410m = cdxi5314m&cdxi5158m;
wire cdxi7411m = cdxi5314m&cdxi5159m;
wire cdxi7412m = cdxi5314m&cdxi5160m;
wire cdxi7413m = cdxi5136m&cdxi5437m;
wire cdxi7414m = cdxi5675m&r30m;
wire cdxi7415m = cdxi5640m&r31m;
wire cdxi7416m = cdxi5083m&cdxi5546m;
wire cdxi7417m = cdxi5533m&r34m;
wire cdxi7418m = cdxi5883m&r35m;
wire cdxi7419m = cdxi5497m&r36m;
wire cdxi7420m = cdxi5424m&r40m;
wire cdxi7421m = cdxi5387m&r41m;
wire cdxi7422m = cdxi5349m&r42m;
wire cdxi7423m = cdxi5534m&r44m;
wire cdxi7424m = cdxi5641m&r45m;
wire cdxi7425m = cdxi5498m&r46m;
wire cdxi7426m = cdxi5425m&r50m;
wire cdxi7427m = cdxi5388m&r51m;
wire cdxi7428m = cdxi5350m&r52m;
wire cdxi7429m = cdxi5426m&r56m;
wire cdxi7430m = cdxi5389m&r57m;
wire cdxi7431m = cdxi5351m&r58m;
wire cdxi7432m = cdxi5314m&r62m;
wire cdxi7433m = cdxi5154m&r64m;
wire cdxi7434m = cdxi4991m&r65m;
wire cdxi7435m = cdxi5136m&r66m;
wire cdxi7436m = cdxi4934m&r70m;
wire cdxi7437m = cdxi5101m&r71m;
wire cdxi7438m = cdxi5083m&r72m;
wire cdxi7439m = cdxi5065m&r76m;
wire cdxi7440m = cdxi4895m&r77m;
wire cdxi7441m = cdxi5028m&r78m;
wire cdxi7442m = cdxi4873m&r82m;
wire cdxi7443m = cdxi4935m&r86m;
wire cdxi7444m = cdxi4896m&r87m;
wire cdxi7445m = cdxi4954m&r88m;
wire cdxi7446m = cdxi4874m&r92m;
wire cdxi7447m = cdxi4875m&r96m;
wire cdxi7448m = cdxi4732m&r101m;
wire cdxi7449m = cdxi4742m&r102m;
wire cdxi7450m = cdxi4762m&r103m;
wire cdxi7451m = cdxi4711m&r107m;
wire cdxi7452m = cdxi4743m&r111m;
wire cdxi7453m = cdxi4712m&r116m;
wire cdxi7454m = (cdxi122m ^ cdxi7392m ^ cdxi7393m ^ cdxi7394m ^ cdxi7395m ^ cdxi7396m ^ cdxi7397m ^ cdxi7398m ^ cdxi7399m ^ cdxi7400m ^ cdxi7401m ^ cdxi7402m ^ cdxi7403m ^ cdxi7404m ^ cdxi7405m ^ cdxi7406m ^ cdxi7407m ^ cdxi7408m ^ cdxi7409m ^ cdxi7410m ^ cdxi7411m ^ cdxi7412m ^ cdxi7413m ^ cdxi7414m ^ cdxi7415m ^ cdxi7416m ^ cdxi7417m ^ cdxi7418m ^ cdxi7419m ^ cdxi7420m ^ cdxi7421m ^ cdxi7422m ^ cdxi7423m ^ cdxi7424m ^ cdxi7425m ^ cdxi7426m ^ cdxi7427m ^ cdxi7428m ^ cdxi7429m ^ cdxi7430m ^ cdxi7431m ^ cdxi7432m ^ cdxi7433m ^ cdxi7434m ^ cdxi7435m ^ cdxi7436m ^ cdxi7437m ^ cdxi7438m ^ cdxi7439m ^ cdxi7440m ^ cdxi7441m ^ cdxi7442m ^ cdxi7443m ^ cdxi7444m ^ cdxi7445m ^ cdxi7446m ^ cdxi7447m ^ cdxi7448m ^ cdxi7449m ^ cdxi7450m ^ cdxi7451m ^ cdxi7452m ^ cdxi7453m);
wire cdxi7455m = a1&cdxi7454m;
wire cdxi7456m = (reg_1_119);
wire cdxi7457m = (reg_1_130);
wire cdxi7458m = reg_1_2&reg_1_3&reg_1_5&reg_1_6&cdxi4738m;
wire cdxi7459m = reg_1_1&cdxi7214m;
wire cdxi7460m = reg_1_1&cdxi7215m;
wire cdxi7461m = reg_1_1&cdxi7216m;
wire cdxi7462m = reg_1_1&cdxi7217m;
wire cdxi7463m = reg_1_1&cdxi7218m;
wire cdxi7464m = reg_1_3&cdxi6685m;
wire cdxi7465m = reg_1_2&reg_1_5&cdxi5698m;
wire cdxi7466m = reg_1_2&reg_1_3&reg_1_6&cdxi5004m;
wire cdxi7467m = reg_1_2&reg_1_3&reg_1_5&reg_1_7&cdxi4905m;
wire cdxi7468m = reg_1_2&reg_1_3&reg_1_5&reg_1_6&cdxi4737m;
wire cdxi7469m = reg_1_1&cdxi7219m;
wire cdxi7470m = reg_1_1&cdxi7220m;
wire cdxi7471m = reg_1_1&cdxi7221m;
wire cdxi7472m = reg_1_1&cdxi7222m;
wire cdxi7473m = reg_1_1&cdxi7223m;
wire cdxi7474m = reg_1_1&cdxi7224m;
wire cdxi7475m = reg_1_1&cdxi7225m;
wire cdxi7476m = reg_1_1&cdxi7226m;
wire cdxi7477m = reg_1_1&cdxi7227m;
wire cdxi7478m = reg_1_1&cdxi7228m;
wire cdxi7479m = reg_1_5&reg_1_6&cdxi5456m;
wire cdxi7480m = reg_1_3&cdxi6695m;
wire cdxi7481m = reg_1_3&cdxi6696m;
wire cdxi7482m = reg_1_3&cdxi6697m;
wire cdxi7483m = reg_1_2&reg_1_6&cdxi5669m;
wire cdxi7484m = reg_1_2&reg_1_5&cdxi5704m;
wire cdxi7485m = reg_1_2&reg_1_5&cdxi5705m;
wire cdxi7486m = reg_1_2&reg_1_3&reg_1_7&cdxi5515m;
wire cdxi7487m = reg_1_2&reg_1_3&reg_1_6&cdxi5000m;
wire cdxi7488m = reg_1_2&reg_1_3&reg_1_5&cdxi5551m;
wire cdxi7489m = reg_1_1&cdxi7229m;
wire cdxi7490m = reg_1_1&cdxi7230m;
wire cdxi7491m = reg_1_1&cdxi7231m;
wire cdxi7492m = reg_1_1&cdxi7232m;
wire cdxi7493m = reg_1_1&cdxi7233m;
wire cdxi7494m = reg_1_1&cdxi7234m;
wire cdxi7495m = reg_1_1&cdxi7235m;
wire cdxi7496m = reg_1_1&cdxi7236m;
wire cdxi7497m = reg_1_1&cdxi7237m;
wire cdxi7498m = reg_1_1&cdxi7238m;
wire cdxi7499m = reg_1_6&cdxi6497m;
wire cdxi7500m = reg_1_5&reg_1_7&cdxi5407m;
wire cdxi7501m = reg_1_5&reg_1_6&cdxi5445m;
wire cdxi7502m = reg_1_3&cdxi6705m;
wire cdxi7503m = reg_1_3&cdxi6706m;
wire cdxi7504m = reg_1_3&cdxi6707m;
wire cdxi7505m = reg_1_2&reg_1_7&cdxi6400m;
wire cdxi7506m = reg_1_2&reg_1_6&cdxi5658m;
wire cdxi7507m = reg_1_2&reg_1_5&cdxi5693m;
wire cdxi7508m = reg_1_2&reg_1_3&cdxi6677m;
wire cdxi7509m = reg_1_1&cdxi7239m;
wire cdxi7510m = reg_1_1&cdxi7240m;
wire cdxi7511m = reg_1_1&cdxi7241m;
wire cdxi7512m = reg_1_1&cdxi7242m;
wire cdxi7513m = reg_1_1&cdxi7243m;
wire cdxi7514m = reg_1_7&cdxi6401m;
wire cdxi7515m = reg_1_6&cdxi6471m;
wire cdxi7516m = reg_1_5&cdxi7320m;
wire cdxi7517m = reg_1_3&cdxi6679m;
wire cdxi7518m = reg_1_2&cdxi7456m;
wire cdxi7519m = reg_1_1&cdxi7213m;
wire cdxi7520m = (cdxi7458m ^ cdxi7459m ^ cdxi7460m ^ cdxi7461m ^ cdxi7462m ^ cdxi7463m ^ cdxi7464m ^ cdxi7465m ^ cdxi7466m ^ cdxi7467m ^ cdxi7468m ^ cdxi7469m ^ cdxi7470m ^ cdxi7471m ^ cdxi7472m ^ cdxi7473m ^ cdxi7474m ^ cdxi7475m ^ cdxi7476m ^ cdxi7477m ^ cdxi7478m ^ cdxi7479m ^ cdxi7480m ^ cdxi7481m ^ cdxi7482m ^ cdxi7483m ^ cdxi7484m ^ cdxi7485m ^ cdxi7486m ^ cdxi7487m ^ cdxi7488m ^ cdxi7489m ^ cdxi7490m ^ cdxi7491m ^ cdxi7492m ^ cdxi7493m ^ cdxi7494m ^ cdxi7495m ^ cdxi7496m ^ cdxi7497m ^ cdxi7498m ^ cdxi7499m ^ cdxi7500m ^ cdxi7501m ^ cdxi7502m ^ cdxi7503m ^ cdxi7504m ^ cdxi7505m ^ cdxi7506m ^ cdxi7507m ^ cdxi7508m ^ cdxi7509m ^ cdxi7510m ^ cdxi7511m ^ cdxi7512m ^ cdxi7513m ^ cdxi7514m ^ cdxi7515m ^ cdxi7516m ^ cdxi7517m ^ cdxi7518m ^ cdxi7519m ^ cdxi7457m);
wire cdxi7521m = reg_1_0&cdxi7520m;
wire cdxi7522m = cdxi5780m&cdxi5154m;
wire cdxi7523m = cdxi4916m&cdxi6017m;
wire cdxi7524m = cdxi4875m&cdxi5710m;
wire cdxi7525m = cdxi4875m&cdxi5950m;
wire cdxi7526m = cdxi6504m&cdxi4733m;
wire cdxi7527m = cdxi6505m&cdxi4790m;
wire cdxi7528m = cdxi4875m&cdxi6191m;
wire cdxi7529m = cdxi4875m&cdxi6192m;
wire cdxi7530m = cdxi4875m&cdxi6193m;
wire cdxi7531m = cdxi4875m&cdxi6194m;
wire cdxi7532m = cdxi4953m&cdxi5539m;
wire cdxi7533m = cdxi5028m&cdxi5750m;
wire cdxi7534m = cdxi5462m&cdxi4995m;
wire cdxi7535m = cdxi4743m&cdxi6854m;
wire cdxi7536m = cdxi6504m&r12m;
wire cdxi7537m = cdxi5498m&cdxi5069m;
wire cdxi7538m = cdxi6573m&r15m;
wire cdxi7539m = cdxi6779m&r16m;
wire cdxi7540m = cdxi6505m&r17m;
wire cdxi7541m = cdxi4875m&cdxi6195m;
wire cdxi7542m = cdxi4875m&cdxi6196m;
wire cdxi7543m = cdxi4875m&cdxi6197m;
wire cdxi7544m = cdxi4875m&cdxi6198m;
wire cdxi7545m = cdxi4875m&cdxi6199m;
wire cdxi7546m = cdxi4875m&cdxi6200m;
wire cdxi7547m = cdxi6017m&r29m;
wire cdxi7548m = cdxi5745m&r30m;
wire cdxi7549m = cdxi4953m&cdxi5545m;
wire cdxi7550m = cdxi4953m&cdxi5546m;
wire cdxi7551m = cdxi5533m&r37m;
wire cdxi7552m = cdxi5883m&r38m;
wire cdxi7553m = cdxi5497m&r39m;
wire cdxi7554m = cdxi5814m&r40m;
wire cdxi7555m = cdxi5462m&r41m;
wire cdxi7556m = cdxi5780m&r42m;
wire cdxi7557m = cdxi5534m&r47m;
wire cdxi7558m = cdxi5641m&r48m;
wire cdxi7559m = cdxi5498m&r49m;
wire cdxi7560m = cdxi5605m&r50m;
wire cdxi7561m = cdxi5463m&r51m;
wire cdxi7562m = cdxi5711m&r52m;
wire cdxi7563m = cdxi5426m&r59m;
wire cdxi7564m = cdxi5389m&r60m;
wire cdxi7565m = cdxi5351m&r61m;
wire cdxi7566m = cdxi5313m&r62m;
wire cdxi7567m = cdxi5154m&r67m;
wire cdxi7568m = cdxi4991m&r68m;
wire cdxi7569m = cdxi5136m&r69m;
wire cdxi7570m = cdxi5064m&r70m;
wire cdxi7571m = cdxi4973m&r71m;
wire cdxi7572m = cdxi4953m&r72m;
wire cdxi7573m = cdxi5065m&r79m;
wire cdxi7574m = cdxi4895m&r80m;
wire cdxi7575m = cdxi5028m&r81m;
wire cdxi7576m = cdxi5009m&r82m;
wire cdxi7577m = cdxi4935m&r89m;
wire cdxi7578m = cdxi4896m&r90m;
wire cdxi7579m = cdxi4954m&r91m;
wire cdxi7580m = cdxi4916m&r92m;
wire cdxi7581m = cdxi4875m&r97m;
wire cdxi7582m = cdxi4732m&r104m;
wire cdxi7583m = cdxi4742m&r105m;
wire cdxi7584m = cdxi4762m&r106m;
wire cdxi7585m = cdxi4722m&r107m;
wire cdxi7586m = cdxi4743m&r112m;
wire cdxi7587m = cdxi4712m&r117m;
wire cdxi7588m = (cdxi123m ^ cdxi7526m ^ cdxi7527m ^ cdxi7528m ^ cdxi7529m ^ cdxi7530m ^ cdxi7531m ^ cdxi7532m ^ cdxi7533m ^ cdxi7534m ^ cdxi7535m ^ cdxi7536m ^ cdxi7537m ^ cdxi7538m ^ cdxi7539m ^ cdxi7540m ^ cdxi7541m ^ cdxi7542m ^ cdxi7543m ^ cdxi7544m ^ cdxi7545m ^ cdxi7546m ^ cdxi7547m ^ cdxi7548m ^ cdxi7549m ^ cdxi7550m ^ cdxi7551m ^ cdxi7552m ^ cdxi7553m ^ cdxi7554m ^ cdxi7555m ^ cdxi7556m ^ cdxi7557m ^ cdxi7558m ^ cdxi7559m ^ cdxi7560m ^ cdxi7561m ^ cdxi7562m ^ cdxi7563m ^ cdxi7564m ^ cdxi7565m ^ cdxi7566m ^ cdxi7567m ^ cdxi7568m ^ cdxi7569m ^ cdxi7570m ^ cdxi7571m ^ cdxi7572m ^ cdxi7573m ^ cdxi7574m ^ cdxi7575m ^ cdxi7576m ^ cdxi7577m ^ cdxi7578m ^ cdxi7579m ^ cdxi7580m ^ cdxi7581m ^ cdxi7582m ^ cdxi7583m ^ cdxi7584m ^ cdxi7585m ^ cdxi7586m ^ cdxi7587m);
wire cdxi7589m = a1&cdxi7588m;
wire cdxi7590m = (reg_1_113);
wire cdxi7591m = (reg_1_131);
wire cdxi7592m = reg_1_2&cdxi6880m;
wire cdxi7593m = reg_1_1&cdxi7079m;
wire cdxi7594m = reg_1_1&cdxi7080m;
wire cdxi7595m = reg_1_1&cdxi7081m;
wire cdxi7596m = reg_1_1&cdxi7082m;
wire cdxi7597m = reg_1_1&cdxi7083m;
wire cdxi7598m = reg_1_4&cdxi6685m;
wire cdxi7599m = reg_1_2&cdxi6885m;
wire cdxi7600m = reg_1_2&cdxi6886m;
wire cdxi7601m = reg_1_2&cdxi6887m;
wire cdxi7602m = reg_1_2&cdxi6888m;
wire cdxi7603m = reg_1_1&cdxi7084m;
wire cdxi7604m = reg_1_1&cdxi7085m;
wire cdxi7605m = reg_1_1&cdxi7086m;
wire cdxi7606m = reg_1_1&cdxi7087m;
wire cdxi7607m = reg_1_1&cdxi7088m;
wire cdxi7608m = reg_1_1&cdxi7089m;
wire cdxi7609m = reg_1_1&cdxi7090m;
wire cdxi7610m = reg_1_1&cdxi7091m;
wire cdxi7611m = reg_1_1&cdxi7092m;
wire cdxi7612m = reg_1_1&cdxi7093m;
wire cdxi7613m = reg_1_5&cdxi6626m;
wire cdxi7614m = reg_1_4&cdxi6695m;
wire cdxi7615m = reg_1_4&cdxi6696m;
wire cdxi7616m = reg_1_4&cdxi6697m;
wire cdxi7617m = reg_1_2&cdxi6895m;
wire cdxi7618m = reg_1_2&cdxi6896m;
wire cdxi7619m = reg_1_2&cdxi6897m;
wire cdxi7620m = reg_1_2&cdxi6898m;
wire cdxi7621m = reg_1_2&cdxi6899m;
wire cdxi7622m = reg_1_2&cdxi6900m;
wire cdxi7623m = reg_1_1&cdxi7094m;
wire cdxi7624m = reg_1_1&cdxi7095m;
wire cdxi7625m = reg_1_1&cdxi7096m;
wire cdxi7626m = reg_1_1&cdxi7097m;
wire cdxi7627m = reg_1_1&cdxi7098m;
wire cdxi7628m = reg_1_1&cdxi7099m;
wire cdxi7629m = reg_1_1&cdxi7100m;
wire cdxi7630m = reg_1_1&cdxi7101m;
wire cdxi7631m = reg_1_1&cdxi7102m;
wire cdxi7632m = reg_1_1&cdxi7103m;
wire cdxi7633m = reg_1_6&reg_1_7&cdxi6261m;
wire cdxi7634m = reg_1_5&cdxi6636m;
wire cdxi7635m = reg_1_5&cdxi6637m;
wire cdxi7636m = reg_1_4&cdxi6705m;
wire cdxi7637m = reg_1_4&cdxi6706m;
wire cdxi7638m = reg_1_4&cdxi6707m;
wire cdxi7639m = reg_1_2&cdxi6905m;
wire cdxi7640m = reg_1_2&cdxi6906m;
wire cdxi7641m = reg_1_2&cdxi6907m;
wire cdxi7642m = reg_1_2&cdxi6908m;
wire cdxi7643m = reg_1_1&cdxi7104m;
wire cdxi7644m = reg_1_1&cdxi7105m;
wire cdxi7645m = reg_1_1&cdxi7106m;
wire cdxi7646m = reg_1_1&cdxi7107m;
wire cdxi7647m = reg_1_1&cdxi7108m;
wire cdxi7648m = reg_1_7&cdxi6539m;
wire cdxi7649m = reg_1_6&cdxi7590m;
wire cdxi7650m = reg_1_5&cdxi6610m;
wire cdxi7651m = reg_1_4&cdxi6679m;
wire cdxi7652m = reg_1_2&cdxi6879m;
wire cdxi7653m = reg_1_1&cdxi7078m;
wire cdxi7654m = (cdxi7592m ^ cdxi7593m ^ cdxi7594m ^ cdxi7595m ^ cdxi7596m ^ cdxi7597m ^ cdxi7598m ^ cdxi7599m ^ cdxi7600m ^ cdxi7601m ^ cdxi7602m ^ cdxi7603m ^ cdxi7604m ^ cdxi7605m ^ cdxi7606m ^ cdxi7607m ^ cdxi7608m ^ cdxi7609m ^ cdxi7610m ^ cdxi7611m ^ cdxi7612m ^ cdxi7613m ^ cdxi7614m ^ cdxi7615m ^ cdxi7616m ^ cdxi7617m ^ cdxi7618m ^ cdxi7619m ^ cdxi7620m ^ cdxi7621m ^ cdxi7622m ^ cdxi7623m ^ cdxi7624m ^ cdxi7625m ^ cdxi7626m ^ cdxi7627m ^ cdxi7628m ^ cdxi7629m ^ cdxi7630m ^ cdxi7631m ^ cdxi7632m ^ cdxi7633m ^ cdxi7634m ^ cdxi7635m ^ cdxi7636m ^ cdxi7637m ^ cdxi7638m ^ cdxi7639m ^ cdxi7640m ^ cdxi7641m ^ cdxi7642m ^ cdxi7643m ^ cdxi7644m ^ cdxi7645m ^ cdxi7646m ^ cdxi7647m ^ cdxi7648m ^ cdxi7649m ^ cdxi7650m ^ cdxi7651m ^ cdxi7652m ^ cdxi7653m ^ cdxi7591m);
wire cdxi7655m = reg_1_0&cdxi7654m;
wire cdxi7656m = cdxi4915m&cdxi6017m;
wire cdxi7657m = cdxi4874m&cdxi5710m;
wire cdxi7658m = cdxi4874m&cdxi5950m;
wire cdxi7659m = cdxi6712m&cdxi4733m;
wire cdxi7660m = cdxi4916m&cdxi6018m;
wire cdxi7661m = cdxi4874m&cdxi6191m;
wire cdxi7662m = cdxi4874m&cdxi6192m;
wire cdxi7663m = cdxi4874m&cdxi6193m;
wire cdxi7664m = cdxi4874m&cdxi6194m;
wire cdxi7665m = cdxi4953m&cdxi5680m;
wire cdxi7666m = cdxi5083m&cdxi5750m;
wire cdxi7667m = cdxi5570m&cdxi4995m;
wire cdxi7668m = cdxi6778m&r11m;
wire cdxi7669m = cdxi6712m&r12m;
wire cdxi7670m = cdxi4954m&cdxi6123m;
wire cdxi7671m = cdxi5463m&cdxi5122m;
wire cdxi7672m = cdxi4916m&cdxi6023m;
wire cdxi7673m = cdxi4916m&cdxi6024m;
wire cdxi7674m = cdxi4874m&cdxi6195m;
wire cdxi7675m = cdxi4874m&cdxi6196m;
wire cdxi7676m = cdxi4874m&cdxi6197m;
wire cdxi7677m = cdxi4874m&cdxi6198m;
wire cdxi7678m = cdxi4874m&cdxi6199m;
wire cdxi7679m = cdxi4874m&cdxi6200m;
wire cdxi7680m = cdxi5136m&cdxi5616m;
wire cdxi7681m = cdxi4973m&cdxi5652m;
wire cdxi7682m = cdxi4953m&cdxi5686m;
wire cdxi7683m = cdxi4953m&cdxi5687m;
wire cdxi7684m = cdxi5675m&r37m;
wire cdxi7685m = cdxi5640m&r38m;
wire cdxi7686m = cdxi5083m&cdxi5757m;
wire cdxi7687m = cdxi5604m&r40m;
wire cdxi7688m = cdxi5570m&r41m;
wire cdxi7689m = cdxi5779m&r42m;
wire cdxi7690m = cdxi5534m&r53m;
wire cdxi7691m = cdxi5641m&r54m;
wire cdxi7692m = cdxi5498m&r55m;
wire cdxi7693m = cdxi5605m&r56m;
wire cdxi7694m = cdxi5463m&r57m;
wire cdxi7695m = cdxi5711m&r58m;
wire cdxi7696m = cdxi5425m&r59m;
wire cdxi7697m = cdxi5388m&r60m;
wire cdxi7698m = cdxi5350m&r61m;
wire cdxi7699m = cdxi5312m&r62m;
wire cdxi7700m = cdxi5154m&r73m;
wire cdxi7701m = cdxi4991m&r74m;
wire cdxi7702m = cdxi5136m&r75m;
wire cdxi7703m = cdxi5064m&r76m;
wire cdxi7704m = cdxi4973m&r77m;
wire cdxi7705m = cdxi4953m&r78m;
wire cdxi7706m = cdxi4934m&r79m;
wire cdxi7707m = cdxi5101m&r80m;
wire cdxi7708m = cdxi5083m&r81m;
wire cdxi7709m = cdxi4915m&r82m;
wire cdxi7710m = cdxi4935m&r93m;
wire cdxi7711m = cdxi4896m&r94m;
wire cdxi7712m = cdxi4954m&r95m;
wire cdxi7713m = cdxi4916m&r96m;
wire cdxi7714m = cdxi4874m&r97m;
wire cdxi7715m = cdxi4732m&r108m;
wire cdxi7716m = cdxi4742m&r109m;
wire cdxi7717m = cdxi4762m&r110m;
wire cdxi7718m = cdxi4722m&r111m;
wire cdxi7719m = cdxi4711m&r112m;
wire cdxi7720m = cdxi4712m&r118m;
wire cdxi7721m = (cdxi124m ^ cdxi7659m ^ cdxi7660m ^ cdxi7661m ^ cdxi7662m ^ cdxi7663m ^ cdxi7664m ^ cdxi7665m ^ cdxi7666m ^ cdxi7667m ^ cdxi7668m ^ cdxi7669m ^ cdxi7670m ^ cdxi7671m ^ cdxi7672m ^ cdxi7673m ^ cdxi7674m ^ cdxi7675m ^ cdxi7676m ^ cdxi7677m ^ cdxi7678m ^ cdxi7679m ^ cdxi7680m ^ cdxi7681m ^ cdxi7682m ^ cdxi7683m ^ cdxi7684m ^ cdxi7685m ^ cdxi7686m ^ cdxi7687m ^ cdxi7688m ^ cdxi7689m ^ cdxi7690m ^ cdxi7691m ^ cdxi7692m ^ cdxi7693m ^ cdxi7694m ^ cdxi7695m ^ cdxi7696m ^ cdxi7697m ^ cdxi7698m ^ cdxi7699m ^ cdxi7700m ^ cdxi7701m ^ cdxi7702m ^ cdxi7703m ^ cdxi7704m ^ cdxi7705m ^ cdxi7706m ^ cdxi7707m ^ cdxi7708m ^ cdxi7709m ^ cdxi7710m ^ cdxi7711m ^ cdxi7712m ^ cdxi7713m ^ cdxi7714m ^ cdxi7715m ^ cdxi7716m ^ cdxi7717m ^ cdxi7718m ^ cdxi7719m ^ cdxi7720m);
wire cdxi7722m = a1&cdxi7721m;
wire cdxi7723m = (reg_1_132);
wire cdxi7724m = reg_1_3&cdxi6880m;
wire cdxi7725m = reg_1_1&cdxi7145m;
wire cdxi7726m = reg_1_1&cdxi7146m;
wire cdxi7727m = reg_1_1&cdxi7147m;
wire cdxi7728m = reg_1_1&cdxi7148m;
wire cdxi7729m = reg_1_1&cdxi7149m;
wire cdxi7730m = reg_1_4&reg_1_5&cdxi5698m;
wire cdxi7731m = reg_1_3&cdxi6885m;
wire cdxi7732m = reg_1_3&cdxi6886m;
wire cdxi7733m = reg_1_3&cdxi6887m;
wire cdxi7734m = reg_1_3&cdxi6888m;
wire cdxi7735m = reg_1_1&cdxi7150m;
wire cdxi7736m = reg_1_1&cdxi7151m;
wire cdxi7737m = reg_1_1&cdxi7152m;
wire cdxi7738m = reg_1_1&cdxi7153m;
wire cdxi7739m = reg_1_1&cdxi7154m;
wire cdxi7740m = reg_1_1&cdxi7155m;
wire cdxi7741m = reg_1_1&cdxi7156m;
wire cdxi7742m = reg_1_1&cdxi7157m;
wire cdxi7743m = reg_1_1&cdxi7158m;
wire cdxi7744m = reg_1_1&cdxi7159m;
wire cdxi7745m = reg_1_5&reg_1_6&cdxi5634m;
wire cdxi7746m = reg_1_4&reg_1_6&cdxi5669m;
wire cdxi7747m = reg_1_4&reg_1_5&cdxi5704m;
wire cdxi7748m = reg_1_4&reg_1_5&cdxi5705m;
wire cdxi7749m = reg_1_3&cdxi6895m;
wire cdxi7750m = reg_1_3&cdxi6896m;
wire cdxi7751m = reg_1_3&cdxi6897m;
wire cdxi7752m = reg_1_3&cdxi6898m;
wire cdxi7753m = reg_1_3&cdxi6899m;
wire cdxi7754m = reg_1_3&cdxi6900m;
wire cdxi7755m = reg_1_1&cdxi7160m;
wire cdxi7756m = reg_1_1&cdxi7161m;
wire cdxi7757m = reg_1_1&cdxi7162m;
wire cdxi7758m = reg_1_1&cdxi7163m;
wire cdxi7759m = reg_1_1&cdxi7164m;
wire cdxi7760m = reg_1_1&cdxi7165m;
wire cdxi7761m = reg_1_1&cdxi7166m;
wire cdxi7762m = reg_1_1&cdxi7167m;
wire cdxi7763m = reg_1_1&cdxi7168m;
wire cdxi7764m = reg_1_1&cdxi7169m;
wire cdxi7765m = reg_1_6&cdxi6839m;
wire cdxi7766m = reg_1_5&reg_1_7&cdxi5587m;
wire cdxi7767m = reg_1_5&reg_1_6&cdxi5623m;
wire cdxi7768m = reg_1_4&reg_1_7&cdxi6400m;
wire cdxi7769m = reg_1_4&reg_1_6&cdxi5658m;
wire cdxi7770m = reg_1_4&reg_1_5&cdxi5693m;
wire cdxi7771m = reg_1_3&cdxi6905m;
wire cdxi7772m = reg_1_3&cdxi6906m;
wire cdxi7773m = reg_1_3&cdxi6907m;
wire cdxi7774m = reg_1_3&cdxi6908m;
wire cdxi7775m = reg_1_1&cdxi7170m;
wire cdxi7776m = reg_1_1&cdxi7171m;
wire cdxi7777m = reg_1_1&cdxi7172m;
wire cdxi7778m = reg_1_1&cdxi7173m;
wire cdxi7779m = reg_1_1&cdxi7174m;
wire cdxi7780m = reg_1_7&cdxi6745m;
wire cdxi7781m = reg_1_6&cdxi6813m;
wire cdxi7782m = reg_1_5&cdxi7321m;
wire cdxi7783m = reg_1_4&cdxi7456m;
wire cdxi7784m = reg_1_3&cdxi6879m;
wire cdxi7785m = reg_1_1&cdxi7144m;
wire cdxi7786m = (cdxi7724m ^ cdxi7725m ^ cdxi7726m ^ cdxi7727m ^ cdxi7728m ^ cdxi7729m ^ cdxi7730m ^ cdxi7731m ^ cdxi7732m ^ cdxi7733m ^ cdxi7734m ^ cdxi7735m ^ cdxi7736m ^ cdxi7737m ^ cdxi7738m ^ cdxi7739m ^ cdxi7740m ^ cdxi7741m ^ cdxi7742m ^ cdxi7743m ^ cdxi7744m ^ cdxi7745m ^ cdxi7746m ^ cdxi7747m ^ cdxi7748m ^ cdxi7749m ^ cdxi7750m ^ cdxi7751m ^ cdxi7752m ^ cdxi7753m ^ cdxi7754m ^ cdxi7755m ^ cdxi7756m ^ cdxi7757m ^ cdxi7758m ^ cdxi7759m ^ cdxi7760m ^ cdxi7761m ^ cdxi7762m ^ cdxi7763m ^ cdxi7764m ^ cdxi7765m ^ cdxi7766m ^ cdxi7767m ^ cdxi7768m ^ cdxi7769m ^ cdxi7770m ^ cdxi7771m ^ cdxi7772m ^ cdxi7773m ^ cdxi7774m ^ cdxi7775m ^ cdxi7776m ^ cdxi7777m ^ cdxi7778m ^ cdxi7779m ^ cdxi7780m ^ cdxi7781m ^ cdxi7782m ^ cdxi7783m ^ cdxi7784m ^ cdxi7785m ^ cdxi7723m);
wire cdxi7787m = reg_1_0&cdxi7786m;
wire cdxi7788m = 0&0 ^ cdxi4743m ^ cdxi4711m ^ cdxi4762m ^ cdxi4732m;
wire cdxi7789m = cdxi4712m&cdxi1m;
wire cdxi7790m = reg_1_1&cdxi4670m;
wire cdxi7791m = cdxi4743m&cdxi2m;
wire cdxi7792m = reg_1_2&cdxi4675m;
wire cdxi7793m = cdxi4743m&cdxi3m;
wire cdxi7794m = reg_1_2&cdxi4680m;
wire cdxi7795m = cdxi4711m&cdxi3m;
wire cdxi7796m = reg_1_3&cdxi4680m;
wire cdxi7797m = cdxi4722m&cdxi4m;
wire cdxi7798m = reg_1_4&cdxi4685m;
wire cdxi7799m = cdxi4762m&cdxi6m;
wire cdxi7800m = reg_1_5&cdxi4699m;
wire cdxi7801m = cdxi4742m&cdxi6m;
wire cdxi7802m = reg_1_6&cdxi4699m;
wire cdxi7803m = cdxi4743m&r0m;
wire cdxi7804m = cdxi4712m&r1m;
wire cdxi7805m = (cdxi7m ^ cdxi7803m ^ cdxi7804m);
wire cdxi7806m = a1&cdxi7805m;
wire cdxi7807m = reg_1_2&cdxi4664m;
wire cdxi7808m = reg_1_1&cdxi4669m;
wire cdxi7809m = (cdxi7807m ^ cdxi7808m ^ cdxi4884m);
wire cdxi7810m = reg_1_0&cdxi7809m;
wire cdxi7811m = cdxi4762m&r0m;
wire cdxi7812m = cdxi4712m&r4m;
wire cdxi7813m = (cdxi10m ^ cdxi7811m ^ cdxi7812m);
wire cdxi7814m = a1&cdxi7813m;
wire cdxi7815m = reg_1_5&cdxi4664m;
wire cdxi7816m = reg_1_1&cdxi4684m;
wire cdxi7817m = (cdxi7815m ^ cdxi7816m ^ cdxi4963m);
wire cdxi7818m = reg_1_0&cdxi7817m;
wire cdxi7819m = cdxi4722m&r1m;
wire cdxi7820m = cdxi4743m&r3m;
wire cdxi7821m = (cdxi14m ^ cdxi7819m ^ cdxi7820m);
wire cdxi7822m = a1&cdxi7821m;
wire cdxi7823m = reg_1_4&cdxi4669m;
wire cdxi7824m = reg_1_2&cdxi4679m;
wire cdxi7825m = (cdxi7823m ^ cdxi7824m ^ cdxi5018m);
wire cdxi7826m = reg_1_0&cdxi7825m;
wire cdxi7827m = cdxi4762m&r1m;
wire cdxi7828m = cdxi4743m&r4m;
wire cdxi7829m = (cdxi15m ^ cdxi7827m ^ cdxi7828m);
wire cdxi7830m = a1&cdxi7829m;
wire cdxi7831m = reg_1_5&cdxi4669m;
wire cdxi7832m = reg_1_2&cdxi4684m;
wire cdxi7833m = (cdxi7831m ^ cdxi7832m ^ cdxi5037m);
wire cdxi7834m = reg_1_0&cdxi7833m;
wire cdxi7835m = a1&cdxi4792m;
wire cdxi7836m = reg_1_0&cdxi4797m;
wire cdxi7837m = a1&cdxi4801m;
wire cdxi7838m = reg_1_0&cdxi4806m;
wire cdxi7839m = a1&cdxi4828m;
wire cdxi7840m = reg_1_0&cdxi4833m;
wire cdxi7841m = a1&cdxi4819m;
wire cdxi7842m = reg_1_0&cdxi4824m;
wire cdxi7843m = a1&cdxi4841m;
wire cdxi7844m = reg_1_0&cdxi4846m;
wire cdxi7845m = a1&cdxi4852m;
wire cdxi7846m = reg_1_0&cdxi4857m;
wire cdxi7847m = cdxi4712m&cdxi7821m;
wire cdxi7848m = reg_1_1&cdxi7825m;
wire cdxi7849m = cdxi4712m&cdxi7829m;
wire cdxi7850m = reg_1_1&cdxi7833m;
wire cdxi7851m = cdxi4712m&cdxi4841m;
wire cdxi7852m = reg_1_1&cdxi4846m;
wire cdxi7853m = cdxi4743m&cdxi4801m;
wire cdxi7854m = reg_1_2&cdxi4806m;
wire cdxi7855m = cdxi4743m&cdxi4810m;
wire cdxi7856m = reg_1_2&cdxi4815m;
wire cdxi7857m = cdxi4743m&cdxi4765m;
wire cdxi7858m = reg_1_2&cdxi4770m;
wire cdxi7859m = cdxi4743m&cdxi4783m;
wire cdxi7860m = reg_1_2&cdxi4788m;
wire cdxi7861m = cdxi4762m&cdxi4852m;
wire cdxi7862m = reg_1_5&cdxi4857m;
wire cdxi7863m = cdxi4743m&cdxi4723m;
wire cdxi7864m = cdxi4916m&r1m;
wire cdxi7865m = cdxi4875m&r3m;
wire cdxi7866m = cdxi4722m&r7m;
wire cdxi7867m = cdxi4743m&r9m;
wire cdxi7868m = cdxi4712m&r14m;
wire cdxi7869m = (cdxi29m ^ cdxi7863m ^ cdxi7864m ^ cdxi7865m ^ cdxi7866m ^ cdxi7867m ^ cdxi7868m);
wire cdxi7870m = a1&cdxi7869m;
wire cdxi7871m = reg_1_2&cdxi4728m;
wire cdxi7872m = reg_1_1&cdxi7823m;
wire cdxi7873m = reg_1_1&cdxi7824m;
wire cdxi7874m = reg_1_4&cdxi4884m;
wire cdxi7875m = reg_1_2&cdxi4727m;
wire cdxi7876m = reg_1_1&cdxi5018m;
wire cdxi7877m = (cdxi7871m ^ cdxi7872m ^ cdxi7873m ^ cdxi7874m ^ cdxi7875m ^ cdxi7876m ^ cdxi5331m);
wire cdxi7878m = reg_1_0&cdxi7877m;
wire cdxi7879m = cdxi4743m&cdxi4733m;
wire cdxi7880m = cdxi4712m&cdxi4790m;
wire cdxi7881m = cdxi4712m&cdxi4791m;
wire cdxi7882m = cdxi4732m&r7m;
wire cdxi7883m = cdxi4743m&r12m;
wire cdxi7884m = cdxi4712m&r17m;
wire cdxi7885m = (cdxi32m ^ cdxi7879m ^ cdxi7880m ^ cdxi7881m ^ cdxi7882m ^ cdxi7883m ^ cdxi7884m);
wire cdxi7886m = a1&cdxi7885m;
wire cdxi7887m = reg_1_2&cdxi4738m;
wire cdxi7888m = reg_1_1&cdxi4795m;
wire cdxi7889m = reg_1_1&cdxi4796m;
wire cdxi7890m = reg_1_7&cdxi4884m;
wire cdxi7891m = reg_1_2&cdxi4737m;
wire cdxi7892m = reg_1_1&cdxi4794m;
wire cdxi7893m = (cdxi7887m ^ cdxi7888m ^ cdxi7889m ^ cdxi7890m ^ cdxi7891m ^ cdxi7892m ^ cdxi5443m);
wire cdxi7894m = reg_1_0&cdxi7893m;
wire cdxi7895m = cdxi5083m&r0m;
wire cdxi7896m = cdxi4712m&cdxi4826m;
wire cdxi7897m = cdxi4712m&cdxi4827m;
wire cdxi7898m = cdxi4762m&r8m;
wire cdxi7899m = cdxi4711m&r10m;
wire cdxi7900m = cdxi4712m&r19m;
wire cdxi7901m = (cdxi34m ^ cdxi7895m ^ cdxi7896m ^ cdxi7897m ^ cdxi7898m ^ cdxi7899m ^ cdxi7900m);
wire cdxi7902m = a1&cdxi7901m;
wire cdxi7903m = reg_1_3&cdxi7815m;
wire cdxi7904m = reg_1_1&cdxi4831m;
wire cdxi7905m = reg_1_1&cdxi4832m;
wire cdxi7906m = reg_1_5&cdxi4717m;
wire cdxi7907m = reg_1_3&cdxi4963m;
wire cdxi7908m = reg_1_1&cdxi4830m;
wire cdxi7909m = (cdxi7903m ^ cdxi7904m ^ cdxi7905m ^ cdxi7906m ^ cdxi7907m ^ cdxi7908m ^ cdxi5369m);
wire cdxi7910m = reg_1_0&cdxi7909m;
wire cdxi7911m = cdxi5101m&r0m;
wire cdxi7912m = cdxi4712m&cdxi4808m;
wire cdxi7913m = cdxi4712m&cdxi4809m;
wire cdxi7914m = cdxi4742m&r8m;
wire cdxi7915m = cdxi4711m&r11m;
wire cdxi7916m = cdxi4712m&r20m;
wire cdxi7917m = (cdxi35m ^ cdxi7911m ^ cdxi7912m ^ cdxi7913m ^ cdxi7914m ^ cdxi7915m ^ cdxi7916m);
wire cdxi7918m = a1&cdxi7917m;
wire cdxi7919m = reg_1_3&reg_1_6&cdxi4664m;
wire cdxi7920m = reg_1_1&cdxi4813m;
wire cdxi7921m = reg_1_1&cdxi4814m;
wire cdxi7922m = reg_1_6&cdxi4717m;
wire cdxi7923m = reg_1_3&cdxi4905m;
wire cdxi7924m = reg_1_1&cdxi4812m;
wire cdxi7925m = (cdxi7919m ^ cdxi7920m ^ cdxi7921m ^ cdxi7922m ^ cdxi7923m ^ cdxi7924m ^ cdxi5406m);
wire cdxi7926m = reg_1_0&cdxi7925m;
wire cdxi7927m = a1&cdxi5195m;
wire cdxi7928m = reg_1_0&cdxi5204m;
wire cdxi7929m = cdxi4711m&cdxi4790m;
wire cdxi7930m = cdxi4743m&cdxi4753m;
wire cdxi7931m = cdxi4743m&cdxi4754m;
wire cdxi7932m = cdxi4732m&r13m;
wire cdxi7933m = cdxi4711m&r17m;
wire cdxi7934m = cdxi4743m&r21m;
wire cdxi7935m = (cdxi46m ^ cdxi7929m ^ cdxi7930m ^ cdxi7931m ^ cdxi7932m ^ cdxi7933m ^ cdxi7934m);
wire cdxi7936m = a1&cdxi7935m;
wire cdxi7937m = reg_1_3&cdxi4795m;
wire cdxi7938m = reg_1_2&cdxi4758m;
wire cdxi7939m = reg_1_2&cdxi4759m;
wire cdxi7940m = reg_1_7&cdxi4885m;
wire cdxi7941m = reg_1_3&cdxi4794m;
wire cdxi7942m = reg_1_2&cdxi4757m;
wire cdxi7943m = (cdxi7937m ^ cdxi7938m ^ cdxi7939m ^ cdxi7940m ^ cdxi7941m ^ cdxi7942m ^ cdxi5444m);
wire cdxi7944m = reg_1_0&cdxi7943m;
wire cdxi7945m = cdxi4742m&cdxi4790m;
wire cdxi7946m = cdxi4743m&cdxi4850m;
wire cdxi7947m = cdxi4743m&cdxi4851m;
wire cdxi7948m = cdxi4732m&r16m;
wire cdxi7949m = cdxi4742m&r17m;
wire cdxi7950m = cdxi4743m&r27m;
wire cdxi7951m = (cdxi52m ^ cdxi7945m ^ cdxi7946m ^ cdxi7947m ^ cdxi7948m ^ cdxi7949m ^ cdxi7950m);
wire cdxi7952m = a1&cdxi7951m;
wire cdxi7953m = reg_1_6&cdxi4795m;
wire cdxi7954m = reg_1_2&cdxi4855m;
wire cdxi7955m = reg_1_2&cdxi4856m;
wire cdxi7956m = reg_1_7&cdxi4748m;
wire cdxi7957m = reg_1_6&cdxi4794m;
wire cdxi7958m = reg_1_2&cdxi4854m;
wire cdxi7959m = (cdxi7953m ^ cdxi7954m ^ cdxi7955m ^ cdxi7956m ^ cdxi7957m ^ cdxi7958m ^ cdxi5552m);
wire cdxi7960m = reg_1_0&cdxi7959m;
wire cdxi7961m = a1&cdxi5275m;
wire cdxi7962m = reg_1_0&cdxi5284m;
wire cdxi7963m = cdxi4762m&cdxi4808m;
wire cdxi7964m = cdxi4711m&cdxi4772m;
wire cdxi7965m = cdxi4711m&cdxi4773m;
wire cdxi7966m = cdxi4742m&r19m;
wire cdxi7967m = cdxi4762m&r20m;
wire cdxi7968m = cdxi4711m&r25m;
wire cdxi7969m = (cdxi56m ^ cdxi7963m ^ cdxi7964m ^ cdxi7965m ^ cdxi7966m ^ cdxi7967m ^ cdxi7968m);
wire cdxi7970m = a1&cdxi7969m;
wire cdxi7971m = reg_1_5&cdxi4813m;
wire cdxi7972m = reg_1_3&cdxi4777m;
wire cdxi7973m = reg_1_3&cdxi4778m;
wire cdxi7974m = reg_1_6&cdxi4830m;
wire cdxi7975m = reg_1_5&cdxi4812m;
wire cdxi7976m = reg_1_3&cdxi4776m;
wire cdxi7977m = (cdxi7971m ^ cdxi7972m ^ cdxi7973m ^ cdxi7974m ^ cdxi7975m ^ cdxi7976m ^ cdxi5865m);
wire cdxi7978m = reg_1_0&cdxi7977m;
wire cdxi7979m = a1&cdxi5298m;
wire cdxi7980m = reg_1_0&cdxi5307m;
wire cdxi7981m = cdxi4712m&cdxi5016m;
wire cdxi7982m = reg_1_1&cdxi5026m;
wire cdxi7983m = cdxi4712m&cdxi7935m;
wire cdxi7984m = reg_1_1&cdxi7943m;
wire cdxi7985m = cdxi4712m&cdxi7951m;
wire cdxi7986m = reg_1_1&cdxi7959m;
wire cdxi7987m = cdxi4712m&cdxi5275m;
wire cdxi7988m = reg_1_1&cdxi5284m;
wire cdxi7989m = cdxi4712m&cdxi7969m;
wire cdxi7990m = reg_1_1&cdxi7977m;
wire cdxi7991m = cdxi4712m&cdxi5161m;
wire cdxi7992m = reg_1_1&cdxi5170m;
wire cdxi7993m = cdxi4743m&cdxi5108m;
wire cdxi7994m = reg_1_2&cdxi5117m;
wire cdxi7995m = cdxi4742m&cdxi4753m;
wire cdxi7996m = cdxi4711m&cdxi4850m;
wire cdxi7997m = cdxi4711m&cdxi4851m;
wire cdxi7998m = cdxi4732m&r20m;
wire cdxi7999m = cdxi4742m&r21m;
wire cdxi8000m = cdxi4711m&r27m;
wire cdxi8001m = (cdxi58m ^ cdxi7995m ^ cdxi7996m ^ cdxi7997m ^ cdxi7998m ^ cdxi7999m ^ cdxi8000m);
wire cdxi8002m = cdxi4743m&cdxi8001m;
wire cdxi8003m = reg_1_6&cdxi4758m;
wire cdxi8004m = reg_1_3&cdxi4855m;
wire cdxi8005m = reg_1_3&cdxi4856m;
wire cdxi8006m = reg_1_7&cdxi4812m;
wire cdxi8007m = reg_1_6&cdxi4757m;
wire cdxi8008m = reg_1_3&cdxi4854m;
wire cdxi8009m = (cdxi8003m ^ cdxi8004m ^ cdxi8005m ^ cdxi8006m ^ cdxi8007m ^ cdxi8008m ^ cdxi5692m);
wire cdxi8010m = reg_1_2&cdxi8009m;
wire cdxi8011m = cdxi4743m&cdxi5298m;
wire cdxi8012m = reg_1_2&cdxi5307m;
wire cdxi8013m = cdxi4711m&cdxi5161m;
wire cdxi8014m = reg_1_3&cdxi5170m;
wire cdxi8015m = cdxi4722m&cdxi5161m;
wire cdxi8016m = reg_1_4&cdxi5170m;
wire cdxi8017m = cdxi5009m&cdxi4733m;
wire cdxi8018m = cdxi4916m&cdxi4790m;
wire cdxi8019m = cdxi4875m&cdxi4839m;
wire cdxi8020m = cdxi4875m&cdxi4840m;
wire cdxi8021m = cdxi5064m&r7m;
wire cdxi8022m = cdxi5065m&r9m;
wire cdxi8023m = cdxi5009m&r12m;
wire cdxi8024m = cdxi4935m&r14m;
wire cdxi8025m = cdxi4916m&r17m;
wire cdxi8026m = cdxi4875m&r24m;
wire cdxi8027m = cdxi4732m&r29m;
wire cdxi8028m = cdxi4722m&r32m;
wire cdxi8029m = cdxi4743m&r39m;
wire cdxi8030m = cdxi4712m&r49m;
wire cdxi8031m = (cdxi69m ^ cdxi8017m ^ cdxi8018m ^ cdxi8019m ^ cdxi8020m ^ cdxi8021m ^ cdxi8022m ^ cdxi8023m ^ cdxi8024m ^ cdxi8025m ^ cdxi8026m ^ cdxi8027m ^ cdxi8028m ^ cdxi8029m ^ cdxi8030m);
wire cdxi8032m = a1&cdxi8031m;
wire cdxi8033m = reg_1_2&reg_1_4&cdxi4738m;
wire cdxi8034m = reg_1_1&cdxi5075m;
wire cdxi8035m = reg_1_1&cdxi5076m;
wire cdxi8036m = reg_1_1&cdxi5077m;
wire cdxi8037m = reg_1_4&cdxi7890m;
wire cdxi8038m = reg_1_2&reg_1_7&cdxi4727m;
wire cdxi8039m = reg_1_2&reg_1_4&cdxi4737m;
wire cdxi8040m = reg_1_1&cdxi5078m;
wire cdxi8041m = reg_1_1&cdxi5079m;
wire cdxi8042m = reg_1_1&cdxi5080m;
wire cdxi8043m = reg_1_7&cdxi5331m;
wire cdxi8044m = reg_1_4&cdxi5443m;
wire cdxi8045m = reg_1_2&cdxi5622m;
wire cdxi8046m = reg_1_1&cdxi5074m;
wire cdxi8047m = (cdxi8033m ^ cdxi8034m ^ cdxi8035m ^ cdxi8036m ^ cdxi8037m ^ cdxi8038m ^ cdxi8039m ^ cdxi8040m ^ cdxi8041m ^ cdxi8042m ^ cdxi8043m ^ cdxi8044m ^ cdxi8045m ^ cdxi8046m ^ cdxi6608m);
wire cdxi8048m = reg_1_0&cdxi8047m;
wire cdxi8049m = cdxi5136m&cdxi4733m;
wire cdxi8050m = cdxi4896m&cdxi4781m;
wire cdxi8051m = cdxi4954m&cdxi4850m;
wire cdxi8052m = cdxi4954m&cdxi4851m;
wire cdxi8053m = cdxi4742m&cdxi4995m;
wire cdxi8054m = cdxi4991m&r11m;
wire cdxi8055m = cdxi5136m&r12m;
wire cdxi8056m = cdxi4935m&r25m;
wire cdxi8057m = cdxi4896m&r26m;
wire cdxi8058m = cdxi4954m&r27m;
wire cdxi8059m = cdxi4732m&r40m;
wire cdxi8060m = cdxi4742m&r41m;
wire cdxi8061m = cdxi4762m&r42m;
wire cdxi8062m = cdxi4712m&r62m;
wire cdxi8063m = (cdxi82m ^ cdxi8049m ^ cdxi8050m ^ cdxi8051m ^ cdxi8052m ^ cdxi8053m ^ cdxi8054m ^ cdxi8055m ^ cdxi8056m ^ cdxi8057m ^ cdxi8058m ^ cdxi8059m ^ cdxi8060m ^ cdxi8061m ^ cdxi8062m);
wire cdxi8064m = a1&cdxi8063m;
wire cdxi8065m = reg_1_5&reg_1_6&cdxi4738m;
wire cdxi8066m = reg_1_1&cdxi5164m;
wire cdxi8067m = reg_1_1&cdxi5165m;
wire cdxi8068m = reg_1_1&cdxi5166m;
wire cdxi8069m = reg_1_6&cdxi5004m;
wire cdxi8070m = reg_1_5&reg_1_7&cdxi4905m;
wire cdxi8071m = reg_1_5&reg_1_6&cdxi4737m;
wire cdxi8072m = reg_1_1&cdxi5167m;
wire cdxi8073m = reg_1_1&cdxi5168m;
wire cdxi8074m = reg_1_1&cdxi5169m;
wire cdxi8075m = reg_1_7&cdxi5515m;
wire cdxi8076m = reg_1_6&cdxi5000m;
wire cdxi8077m = reg_1_5&cdxi5551m;
wire cdxi8078m = reg_1_1&cdxi5163m;
wire cdxi8079m = (cdxi8065m ^ cdxi8066m ^ cdxi8067m ^ cdxi8068m ^ cdxi8069m ^ cdxi8070m ^ cdxi8071m ^ cdxi8072m ^ cdxi8073m ^ cdxi8074m ^ cdxi8075m ^ cdxi8076m ^ cdxi8077m ^ cdxi8078m ^ cdxi6677m);
wire cdxi8080m = reg_1_0&cdxi8079m;
wire cdxi8081m = cdxi4973m&cdxi4790m;
wire cdxi8082m = cdxi4895m&cdxi4839m;
wire cdxi8083m = cdxi5009m&cdxi4850m;
wire cdxi8084m = cdxi5009m&cdxi4851m;
wire cdxi8085m = cdxi4742m&cdxi5069m;
wire cdxi8086m = cdxi5064m&r16m;
wire cdxi8087m = cdxi4973m&r17m;
wire cdxi8088m = cdxi5065m&r23m;
wire cdxi8089m = cdxi4895m&r24m;
wire cdxi8090m = cdxi5009m&r27m;
wire cdxi8091m = cdxi4732m&r48m;
wire cdxi8092m = cdxi4742m&r49m;
wire cdxi8093m = cdxi4722m&r52m;
wire cdxi8094m = cdxi4743m&r61m;
wire cdxi8095m = (cdxi91m ^ cdxi8081m ^ cdxi8082m ^ cdxi8083m ^ cdxi8084m ^ cdxi8085m ^ cdxi8086m ^ cdxi8087m ^ cdxi8088m ^ cdxi8089m ^ cdxi8090m ^ cdxi8091m ^ cdxi8092m ^ cdxi8093m ^ cdxi8094m);
wire cdxi8096m = a1&cdxi8095m;
wire cdxi8097m = reg_1_4&cdxi7953m;
wire cdxi8098m = reg_1_2&cdxi5259m;
wire cdxi8099m = reg_1_2&cdxi5260m;
wire cdxi8100m = reg_1_2&cdxi5261m;
wire cdxi8101m = reg_1_6&cdxi5078m;
wire cdxi8102m = reg_1_4&cdxi7956m;
wire cdxi8103m = reg_1_4&cdxi7957m;
wire cdxi8104m = reg_1_2&cdxi5262m;
wire cdxi8105m = reg_1_2&cdxi5263m;
wire cdxi8106m = reg_1_2&cdxi5264m;
wire cdxi8107m = reg_1_7&cdxi5055m;
wire cdxi8108m = reg_1_6&cdxi5074m;
wire cdxi8109m = reg_1_4&cdxi5552m;
wire cdxi8110m = reg_1_2&cdxi5258m;
wire cdxi8111m = (cdxi8097m ^ cdxi8098m ^ cdxi8099m ^ cdxi8100m ^ cdxi8101m ^ cdxi8102m ^ cdxi8103m ^ cdxi8104m ^ cdxi8105m ^ cdxi8106m ^ cdxi8107m ^ cdxi8108m ^ cdxi8109m ^ cdxi8110m ^ cdxi6609m);
wire cdxi8112m = reg_1_0&cdxi8111m;
wire cdxi8113m = cdxi5136m&cdxi4790m;
wire cdxi8114m = cdxi4895m&cdxi4781m;
wire cdxi8115m = cdxi5028m&cdxi4850m;
wire cdxi8116m = cdxi5028m&cdxi4851m;
wire cdxi8117m = cdxi5154m&r15m;
wire cdxi8118m = cdxi4991m&r16m;
wire cdxi8119m = cdxi5136m&r17m;
wire cdxi8120m = cdxi5065m&r25m;
wire cdxi8121m = cdxi4895m&r26m;
wire cdxi8122m = cdxi5028m&r27m;
wire cdxi8123m = cdxi4732m&r50m;
wire cdxi8124m = cdxi4742m&r51m;
wire cdxi8125m = cdxi4762m&r52m;
wire cdxi8126m = cdxi4743m&r62m;
wire cdxi8127m = (cdxi92m ^ cdxi8113m ^ cdxi8114m ^ cdxi8115m ^ cdxi8116m ^ cdxi8117m ^ cdxi8118m ^ cdxi8119m ^ cdxi8120m ^ cdxi8121m ^ cdxi8122m ^ cdxi8123m ^ cdxi8124m ^ cdxi8125m ^ cdxi8126m);
wire cdxi8128m = a1&cdxi8127m;
wire cdxi8129m = reg_1_5&cdxi7953m;
wire cdxi8130m = reg_1_2&cdxi5164m;
wire cdxi8131m = reg_1_2&cdxi5165m;
wire cdxi8132m = reg_1_2&cdxi5166m;
wire cdxi8133m = reg_1_6&cdxi5239m;
wire cdxi8134m = reg_1_5&cdxi7956m;
wire cdxi8135m = reg_1_5&cdxi7957m;
wire cdxi8136m = reg_1_2&cdxi5167m;
wire cdxi8137m = reg_1_2&cdxi5168m;
wire cdxi8138m = reg_1_2&cdxi5169m;
wire cdxi8139m = reg_1_7&cdxi5218m;
wire cdxi8140m = reg_1_6&cdxi5235m;
wire cdxi8141m = reg_1_5&cdxi5552m;
wire cdxi8142m = reg_1_2&cdxi5163m;
wire cdxi8143m = (cdxi8129m ^ cdxi8130m ^ cdxi8131m ^ cdxi8132m ^ cdxi8133m ^ cdxi8134m ^ cdxi8135m ^ cdxi8136m ^ cdxi8137m ^ cdxi8138m ^ cdxi8139m ^ cdxi8140m ^ cdxi8141m ^ cdxi8142m ^ cdxi6678m);
wire cdxi8144m = reg_1_0&cdxi8143m;
wire cdxi8145m = a1&cdxi6133m;
wire cdxi8146m = reg_1_0&cdxi6150m;
wire cdxi8147m = a1&cdxi6205m;
wire cdxi8148m = reg_1_0&cdxi6222m;
wire cdxi8149m = cdxi4712m&cdxi5795m;
wire cdxi8150m = reg_1_1&cdxi5812m;
wire cdxi8151m = cdxi4712m&cdxi5863m;
wire cdxi8152m = reg_1_1&cdxi5881m;
wire cdxi8153m = cdxi4712m&cdxi5898m;
wire cdxi8154m = reg_1_1&cdxi5915m;
wire cdxi8155m = cdxi4712m&cdxi8127m;
wire cdxi8156m = reg_1_1&cdxi8143m;
wire cdxi8157m = cdxi4712m&cdxi6032m;
wire cdxi8158m = reg_1_1&cdxi6049m;
wire cdxi8159m = cdxi4712m&cdxi6205m;
wire cdxi8160m = reg_1_1&cdxi6222m;
wire cdxi8161m = cdxi4743m&cdxi6205m;
wire cdxi8162m = reg_1_2&cdxi6222m;
wire cdxi8163m = cdxi5387m&cdxi4733m;
wire cdxi8164m = cdxi5388m&cdxi4790m;
wire cdxi8165m = cdxi5389m&cdxi4753m;
wire cdxi8166m = cdxi5314m&cdxi4850m;
wire cdxi8167m = cdxi5314m&cdxi4851m;
wire cdxi8168m = cdxi5675m&r7m;
wire cdxi8169m = cdxi4895m&cdxi4939m;
wire cdxi8170m = cdxi5424m&r11m;
wire cdxi8171m = cdxi5387m&r12m;
wire cdxi8172m = cdxi5534m&r13m;
wire cdxi8173m = cdxi5425m&r16m;
wire cdxi8174m = cdxi5388m&r17m;
wire cdxi8175m = cdxi5426m&r20m;
wire cdxi8176m = cdxi5389m&r21m;
wire cdxi8177m = cdxi5314m&r27m;
wire cdxi8178m = cdxi5154m&r28m;
wire cdxi8179m = cdxi4934m&r31m;
wire cdxi8180m = cdxi5101m&r32m;
wire cdxi8181m = cdxi5065m&r35m;
wire cdxi8182m = cdxi4895m&r36m;
wire cdxi8183m = cdxi4873m&r42m;
wire cdxi8184m = cdxi4935m&r45m;
wire cdxi8185m = cdxi4896m&r46m;
wire cdxi8186m = cdxi4874m&r52m;
wire cdxi8187m = cdxi4875m&r58m;
wire cdxi8188m = cdxi4732m&r65m;
wire cdxi8189m = cdxi4742m&r66m;
wire cdxi8190m = cdxi4711m&r72m;
wire cdxi8191m = cdxi4743m&r78m;
wire cdxi8192m = cdxi4712m&r88m;
wire cdxi8193m = (cdxi103m ^ cdxi8163m ^ cdxi8164m ^ cdxi8165m ^ cdxi8166m ^ cdxi8167m ^ cdxi8168m ^ cdxi8169m ^ cdxi8170m ^ cdxi8171m ^ cdxi8172m ^ cdxi8173m ^ cdxi8174m ^ cdxi8175m ^ cdxi8176m ^ cdxi8177m ^ cdxi8178m ^ cdxi8179m ^ cdxi8180m ^ cdxi8181m ^ cdxi8182m ^ cdxi8183m ^ cdxi8184m ^ cdxi8185m ^ cdxi8186m ^ cdxi8187m ^ cdxi8188m ^ cdxi8189m ^ cdxi8190m ^ cdxi8191m ^ cdxi8192m);
wire cdxi8194m = a1&cdxi8193m;
wire cdxi8195m = reg_1_2&cdxi5694m;
wire cdxi8196m = reg_1_1&cdxi5934m;
wire cdxi8197m = reg_1_1&cdxi5935m;
wire cdxi8198m = reg_1_1&cdxi5936m;
wire cdxi8199m = reg_1_1&cdxi5937m;
wire cdxi8200m = reg_1_3&cdxi5558m;
wire cdxi8201m = reg_1_2&cdxi5698m;
wire cdxi8202m = reg_1_2&cdxi5699m;
wire cdxi8203m = reg_1_2&cdxi5700m;
wire cdxi8204m = reg_1_1&cdxi5938m;
wire cdxi8205m = reg_1_1&cdxi5939m;
wire cdxi8206m = reg_1_1&cdxi5940m;
wire cdxi8207m = reg_1_1&cdxi5941m;
wire cdxi8208m = reg_1_1&cdxi5942m;
wire cdxi8209m = reg_1_1&cdxi5943m;
wire cdxi8210m = reg_1_6&cdxi5456m;
wire cdxi8211m = reg_1_3&cdxi5564m;
wire cdxi8212m = reg_1_3&cdxi5565m;
wire cdxi8213m = reg_1_2&cdxi5704m;
wire cdxi8214m = reg_1_2&cdxi5705m;
wire cdxi8215m = reg_1_2&cdxi5706m;
wire cdxi8216m = reg_1_1&cdxi5944m;
wire cdxi8217m = reg_1_1&cdxi5945m;
wire cdxi8218m = reg_1_1&cdxi5946m;
wire cdxi8219m = reg_1_1&cdxi5947m;
wire cdxi8220m = reg_1_7&cdxi5407m;
wire cdxi8221m = reg_1_6&cdxi5445m;
wire cdxi8222m = reg_1_3&cdxi5553m;
wire cdxi8223m = reg_1_2&cdxi5693m;
wire cdxi8224m = reg_1_1&cdxi5933m;
wire cdxi8225m = (cdxi8195m ^ cdxi8196m ^ cdxi8197m ^ cdxi8198m ^ cdxi8199m ^ cdxi8200m ^ cdxi8201m ^ cdxi8202m ^ cdxi8203m ^ cdxi8204m ^ cdxi8205m ^ cdxi8206m ^ cdxi8207m ^ cdxi8208m ^ cdxi8209m ^ cdxi8210m ^ cdxi8211m ^ cdxi8212m ^ cdxi8213m ^ cdxi8214m ^ cdxi8215m ^ cdxi8216m ^ cdxi8217m ^ cdxi8218m ^ cdxi8219m ^ cdxi8220m ^ cdxi8221m ^ cdxi8222m ^ cdxi8223m ^ cdxi8224m ^ cdxi7320m);
wire cdxi8226m = reg_1_0&cdxi8225m;
wire cdxi8227m = cdxi4915m&cdxi5210m;
wire cdxi8228m = cdxi5780m&cdxi4808m;
wire cdxi8229m = cdxi4873m&cdxi5137m;
wire cdxi8230m = cdxi4873m&cdxi5138m;
wire cdxi8231m = cdxi4873m&cdxi5139m;
wire cdxi8232m = cdxi4953m&cdxi5192m;
wire cdxi8233m = cdxi5083m&cdxi5050m;
wire cdxi8234m = cdxi4915m&cdxi5213m;
wire cdxi8235m = cdxi4915m&cdxi5214m;
wire cdxi8236m = cdxi5028m&cdxi5105m;
wire cdxi8237m = cdxi5462m&r19m;
wire cdxi8238m = cdxi5780m&r20m;
wire cdxi8239m = cdxi4873m&cdxi5140m;
wire cdxi8240m = cdxi4873m&cdxi5141m;
wire cdxi8241m = cdxi4873m&cdxi5142m;
wire cdxi8242m = cdxi5136m&r43m;
wire cdxi8243m = cdxi4973m&r44m;
wire cdxi8244m = cdxi4953m&r45m;
wire cdxi8245m = cdxi5101m&r47m;
wire cdxi8246m = cdxi5083m&r48m;
wire cdxi8247m = cdxi4915m&r50m;
wire cdxi8248m = cdxi4895m&r53m;
wire cdxi8249m = cdxi5028m&r54m;
wire cdxi8250m = cdxi5009m&r56m;
wire cdxi8251m = cdxi4873m&r59m;
wire cdxi8252m = cdxi4742m&r83m;
wire cdxi8253m = cdxi4762m&r84m;
wire cdxi8254m = cdxi4722m&r86m;
wire cdxi8255m = cdxi4711m&r89m;
wire cdxi8256m = cdxi4743m&r93m;
wire cdxi8257m = (cdxi113m ^ cdxi8227m ^ cdxi8228m ^ cdxi8229m ^ cdxi8230m ^ cdxi8231m ^ cdxi8232m ^ cdxi8233m ^ cdxi8234m ^ cdxi8235m ^ cdxi8236m ^ cdxi8237m ^ cdxi8238m ^ cdxi8239m ^ cdxi8240m ^ cdxi8241m ^ cdxi8242m ^ cdxi8243m ^ cdxi8244m ^ cdxi8245m ^ cdxi8246m ^ cdxi8247m ^ cdxi8248m ^ cdxi8249m ^ cdxi8250m ^ cdxi8251m ^ cdxi8252m ^ cdxi8253m ^ cdxi8254m ^ cdxi8255m ^ cdxi8256m);
wire cdxi8258m = a1&cdxi8257m;
wire cdxi8259m = (reg_1_121);
wire cdxi8260m = reg_1_3&cdxi5968m;
wire cdxi8261m = reg_1_2&cdxi6169m;
wire cdxi8262m = reg_1_2&cdxi6170m;
wire cdxi8263m = reg_1_2&cdxi6171m;
wire cdxi8264m = reg_1_2&cdxi6172m;
wire cdxi8265m = reg_1_4&cdxi5871m;
wire cdxi8266m = reg_1_3&cdxi5972m;
wire cdxi8267m = reg_1_3&cdxi5973m;
wire cdxi8268m = reg_1_3&cdxi5974m;
wire cdxi8269m = reg_1_2&cdxi6173m;
wire cdxi8270m = reg_1_2&cdxi6174m;
wire cdxi8271m = reg_1_2&cdxi6175m;
wire cdxi8272m = reg_1_2&cdxi6176m;
wire cdxi8273m = reg_1_2&cdxi6177m;
wire cdxi8274m = reg_1_2&cdxi6178m;
wire cdxi8275m = reg_1_5&cdxi6078m;
wire cdxi8276m = reg_1_4&cdxi5877m;
wire cdxi8277m = reg_1_4&cdxi5878m;
wire cdxi8278m = reg_1_3&cdxi5978m;
wire cdxi8279m = reg_1_3&cdxi5979m;
wire cdxi8280m = reg_1_3&cdxi5980m;
wire cdxi8281m = reg_1_2&cdxi6179m;
wire cdxi8282m = reg_1_2&cdxi6180m;
wire cdxi8283m = reg_1_2&cdxi6181m;
wire cdxi8284m = reg_1_2&cdxi6182m;
wire cdxi8285m = reg_1_6&cdxi5797m;
wire cdxi8286m = reg_1_5&cdxi6067m;
wire cdxi8287m = reg_1_4&cdxi5866m;
wire cdxi8288m = reg_1_3&cdxi5967m;
wire cdxi8289m = reg_1_2&cdxi6168m;
wire cdxi8290m = (cdxi8260m ^ cdxi8261m ^ cdxi8262m ^ cdxi8263m ^ cdxi8264m ^ cdxi8265m ^ cdxi8266m ^ cdxi8267m ^ cdxi8268m ^ cdxi8269m ^ cdxi8270m ^ cdxi8271m ^ cdxi8272m ^ cdxi8273m ^ cdxi8274m ^ cdxi8275m ^ cdxi8276m ^ cdxi8277m ^ cdxi8278m ^ cdxi8279m ^ cdxi8280m ^ cdxi8281m ^ cdxi8282m ^ cdxi8283m ^ cdxi8284m ^ cdxi8285m ^ cdxi8286m ^ cdxi8287m ^ cdxi8288m ^ cdxi8289m ^ cdxi8259m);
wire cdxi8291m = reg_1_0&cdxi8290m;
wire cdxi8292m = cdxi4873m&cdxi5950m;
wire cdxi8293m = cdxi5314m&cdxi4953m;
wire cdxi8294m = cdxi8292m&r0m;
wire cdxi8295m = cdxi4874m&cdxi5951m;
wire cdxi8296m = cdxi4875m&cdxi6152m;
wire cdxi8297m = cdxi5314m&cdxi5137m;
wire cdxi8298m = cdxi5314m&cdxi5138m;
wire cdxi8299m = cdxi5314m&cdxi5139m;
wire cdxi8300m = cdxi4915m&cdxi5503m;
wire cdxi8301m = cdxi6504m&r8m;
wire cdxi8302m = cdxi5349m&cdxi4977m;
wire cdxi8303m = cdxi6296m&r10m;
wire cdxi8304m = cdxi6224m&r11m;
wire cdxi8305m = cdxi4916m&cdxi5853m;
wire cdxi8306m = cdxi5350m&cdxi5050m;
wire cdxi8307m = cdxi4874m&cdxi5956m;
wire cdxi8308m = cdxi4874m&cdxi5957m;
wire cdxi8309m = cdxi5351m&cdxi5105m;
wire cdxi8310m = cdxi4875m&cdxi6157m;
wire cdxi8311m = cdxi4875m&cdxi6158m;
wire cdxi8312m = cdxi5314m&cdxi5140m;
wire cdxi8313m = cdxi5314m&cdxi5141m;
wire cdxi8314m = cdxi5314m&cdxi5142m;
wire cdxi8315m = cdxi4953m&cdxi5400m;
wire cdxi8316m = cdxi5083m&cdxi5474m;
wire cdxi8317m = cdxi4915m&cdxi5509m;
wire cdxi8318m = cdxi4915m&cdxi5510m;
wire cdxi8319m = cdxi5497m&r33m;
wire cdxi8320m = cdxi5462m&r34m;
wire cdxi8321m = cdxi5780m&r35m;
wire cdxi8322m = cdxi5387m&r37m;
wire cdxi8323m = cdxi5349m&r38m;
wire cdxi8324m = cdxi5311m&r40m;
wire cdxi8325m = cdxi5498m&r43m;
wire cdxi8326m = cdxi5463m&r44m;
wire cdxi8327m = cdxi5711m&r45m;
wire cdxi8328m = cdxi5388m&r47m;
wire cdxi8329m = cdxi5350m&r48m;
wire cdxi8330m = cdxi5312m&r50m;
wire cdxi8331m = cdxi5389m&r53m;
wire cdxi8332m = cdxi5351m&r54m;
wire cdxi8333m = cdxi5313m&r56m;
wire cdxi8334m = cdxi5314m&r59m;
wire cdxi8335m = cdxi5136m&r63m;
wire cdxi8336m = cdxi4973m&r64m;
wire cdxi8337m = cdxi4953m&r65m;
wire cdxi8338m = cdxi5101m&r67m;
wire cdxi8339m = cdxi5083m&r68m;
wire cdxi8340m = cdxi4915m&r70m;
wire cdxi8341m = cdxi4895m&r73m;
wire cdxi8342m = cdxi5028m&r74m;
wire cdxi8343m = cdxi5009m&r76m;
wire cdxi8344m = cdxi4873m&r79m;
wire cdxi8345m = cdxi4896m&r83m;
wire cdxi8346m = cdxi4954m&r84m;
wire cdxi8347m = cdxi4916m&r86m;
wire cdxi8348m = cdxi4874m&r89m;
wire cdxi8349m = cdxi4875m&r93m;
wire cdxi8350m = cdxi4742m&r98m;
wire cdxi8351m = cdxi4762m&r99m;
wire cdxi8352m = cdxi4722m&r101m;
wire cdxi8353m = cdxi4711m&r104m;
wire cdxi8354m = cdxi4743m&r108m;
wire cdxi8355m = cdxi4712m&r113m;
wire cdxi8356m = (cdxi119m ^ cdxi8294m ^ cdxi8295m ^ cdxi8296m ^ cdxi8297m ^ cdxi8298m ^ cdxi8299m ^ cdxi8300m ^ cdxi8301m ^ cdxi8302m ^ cdxi8303m ^ cdxi8304m ^ cdxi8305m ^ cdxi8306m ^ cdxi8307m ^ cdxi8308m ^ cdxi8309m ^ cdxi8310m ^ cdxi8311m ^ cdxi8312m ^ cdxi8313m ^ cdxi8314m ^ cdxi8315m ^ cdxi8316m ^ cdxi8317m ^ cdxi8318m ^ cdxi8319m ^ cdxi8320m ^ cdxi8321m ^ cdxi8322m ^ cdxi8323m ^ cdxi8324m ^ cdxi8325m ^ cdxi8326m ^ cdxi8327m ^ cdxi8328m ^ cdxi8329m ^ cdxi8330m ^ cdxi8331m ^ cdxi8332m ^ cdxi8333m ^ cdxi8334m ^ cdxi8335m ^ cdxi8336m ^ cdxi8337m ^ cdxi8338m ^ cdxi8339m ^ cdxi8340m ^ cdxi8341m ^ cdxi8342m ^ cdxi8343m ^ cdxi8344m ^ cdxi8345m ^ cdxi8346m ^ cdxi8347m ^ cdxi8348m ^ cdxi8349m ^ cdxi8350m ^ cdxi8351m ^ cdxi8352m ^ cdxi8353m ^ cdxi8354m ^ cdxi8355m);
wire cdxi8357m = a1&cdxi8356m;
wire cdxi8358m = (reg_1_127);
wire cdxi8359m = reg_1_2&cdxi6746m;
wire cdxi8360m = reg_1_1&cdxi8260m;
wire cdxi8361m = reg_1_1&cdxi8261m;
wire cdxi8362m = reg_1_1&cdxi8262m;
wire cdxi8363m = reg_1_1&cdxi8263m;
wire cdxi8364m = reg_1_1&cdxi8264m;
wire cdxi8365m = reg_1_3&cdxi6545m;
wire cdxi8366m = reg_1_2&cdxi6751m;
wire cdxi8367m = reg_1_2&cdxi6752m;
wire cdxi8368m = reg_1_2&cdxi6753m;
wire cdxi8369m = reg_1_2&cdxi6754m;
wire cdxi8370m = reg_1_1&cdxi8265m;
wire cdxi8371m = reg_1_1&cdxi8266m;
wire cdxi8372m = reg_1_1&cdxi8267m;
wire cdxi8373m = reg_1_1&cdxi8268m;
wire cdxi8374m = reg_1_1&cdxi8269m;
wire cdxi8375m = reg_1_1&cdxi8270m;
wire cdxi8376m = reg_1_1&cdxi8271m;
wire cdxi8377m = reg_1_1&cdxi8272m;
wire cdxi8378m = reg_1_1&cdxi8273m;
wire cdxi8379m = reg_1_1&cdxi8274m;
wire cdxi8380m = reg_1_4&cdxi6417m;
wire cdxi8381m = reg_1_3&cdxi6555m;
wire cdxi8382m = reg_1_3&cdxi6556m;
wire cdxi8383m = reg_1_3&cdxi6557m;
wire cdxi8384m = reg_1_2&cdxi6761m;
wire cdxi8385m = reg_1_2&cdxi6762m;
wire cdxi8386m = reg_1_2&cdxi6763m;
wire cdxi8387m = reg_1_2&cdxi6764m;
wire cdxi8388m = reg_1_2&cdxi6765m;
wire cdxi8389m = reg_1_2&cdxi6766m;
wire cdxi8390m = reg_1_1&cdxi8275m;
wire cdxi8391m = reg_1_1&cdxi8276m;
wire cdxi8392m = reg_1_1&cdxi8277m;
wire cdxi8393m = reg_1_1&cdxi8278m;
wire cdxi8394m = reg_1_1&cdxi8279m;
wire cdxi8395m = reg_1_1&cdxi8280m;
wire cdxi8396m = reg_1_1&cdxi8281m;
wire cdxi8397m = reg_1_1&cdxi8282m;
wire cdxi8398m = reg_1_1&cdxi8283m;
wire cdxi8399m = reg_1_1&cdxi8284m;
wire cdxi8400m = reg_1_5&cdxi6358m;
wire cdxi8401m = reg_1_4&cdxi6427m;
wire cdxi8402m = reg_1_4&cdxi6428m;
wire cdxi8403m = reg_1_3&cdxi6565m;
wire cdxi8404m = reg_1_3&cdxi6566m;
wire cdxi8405m = reg_1_3&cdxi6567m;
wire cdxi8406m = reg_1_2&cdxi6771m;
wire cdxi8407m = reg_1_2&cdxi6772m;
wire cdxi8408m = reg_1_2&cdxi6773m;
wire cdxi8409m = reg_1_2&cdxi6774m;
wire cdxi8410m = reg_1_1&cdxi8285m;
wire cdxi8411m = reg_1_1&cdxi8286m;
wire cdxi8412m = reg_1_1&cdxi8287m;
wire cdxi8413m = reg_1_1&cdxi8288m;
wire cdxi8414m = reg_1_1&cdxi8289m;
wire cdxi8415m = reg_1_6&cdxi6263m;
wire cdxi8416m = reg_1_5&cdxi6332m;
wire cdxi8417m = reg_1_4&cdxi6401m;
wire cdxi8418m = reg_1_3&cdxi6539m;
wire cdxi8419m = reg_1_2&cdxi6745m;
wire cdxi8420m = reg_1_1&cdxi8259m;
wire cdxi8421m = (cdxi8359m ^ cdxi8360m ^ cdxi8361m ^ cdxi8362m ^ cdxi8363m ^ cdxi8364m ^ cdxi8365m ^ cdxi8366m ^ cdxi8367m ^ cdxi8368m ^ cdxi8369m ^ cdxi8370m ^ cdxi8371m ^ cdxi8372m ^ cdxi8373m ^ cdxi8374m ^ cdxi8375m ^ cdxi8376m ^ cdxi8377m ^ cdxi8378m ^ cdxi8379m ^ cdxi8380m ^ cdxi8381m ^ cdxi8382m ^ cdxi8383m ^ cdxi8384m ^ cdxi8385m ^ cdxi8386m ^ cdxi8387m ^ cdxi8388m ^ cdxi8389m ^ cdxi8390m ^ cdxi8391m ^ cdxi8392m ^ cdxi8393m ^ cdxi8394m ^ cdxi8395m ^ cdxi8396m ^ cdxi8397m ^ cdxi8398m ^ cdxi8399m ^ cdxi8400m ^ cdxi8401m ^ cdxi8402m ^ cdxi8403m ^ cdxi8404m ^ cdxi8405m ^ cdxi8406m ^ cdxi8407m ^ cdxi8408m ^ cdxi8409m ^ cdxi8410m ^ cdxi8411m ^ cdxi8412m ^ cdxi8413m ^ cdxi8414m ^ cdxi8415m ^ cdxi8416m ^ cdxi8417m ^ cdxi8418m ^ cdxi8419m ^ cdxi8420m ^ cdxi8358m);
wire cdxi8422m = reg_1_0&cdxi8421m;
wire cdxi8423m = cdxi4873m&cdxi5710m;
wire cdxi8424m = cdxi6712m&cdxi4790m;
wire cdxi8425m = cdxi6504m&cdxi4753m;
wire cdxi8426m = cdxi4873m&cdxi6191m;
wire cdxi8427m = cdxi4873m&cdxi6192m;
wire cdxi8428m = cdxi4873m&cdxi6193m;
wire cdxi8429m = cdxi4873m&cdxi6194m;
wire cdxi8430m = cdxi4953m&cdxi5921m;
wire cdxi8431m = cdxi5848m&cdxi5069m;
wire cdxi8432m = cdxi6979m&r15m;
wire cdxi8433m = cdxi6778m&r16m;
wire cdxi8434m = cdxi6712m&r17m;
wire cdxi8435m = cdxi5028m&cdxi6123m;
wire cdxi8436m = cdxi5462m&cdxi5122m;
wire cdxi8437m = cdxi6912m&r20m;
wire cdxi8438m = cdxi6504m&r21m;
wire cdxi8439m = cdxi4873m&cdxi6195m;
wire cdxi8440m = cdxi4873m&cdxi6196m;
wire cdxi8441m = cdxi4873m&cdxi6197m;
wire cdxi8442m = cdxi4873m&cdxi6198m;
wire cdxi8443m = cdxi4873m&cdxi6199m;
wire cdxi8444m = cdxi4873m&cdxi6200m;
wire cdxi8445m = cdxi5136m&cdxi5825m;
wire cdxi8446m = cdxi5745m&r44m;
wire cdxi8447m = cdxi5710m&r45m;
wire cdxi8448m = cdxi4953m&cdxi5928m;
wire cdxi8449m = cdxi5675m&r47m;
wire cdxi8450m = cdxi5640m&r48m;
wire cdxi8451m = cdxi5848m&r49m;
wire cdxi8452m = cdxi5604m&r50m;
wire cdxi8453m = cdxi5570m&r51m;
wire cdxi8454m = cdxi5779m&r52m;
wire cdxi8455m = cdxi5533m&r53m;
wire cdxi8456m = cdxi5883m&r54m;
wire cdxi8457m = cdxi5497m&r55m;
wire cdxi8458m = cdxi5814m&r56m;
wire cdxi8459m = cdxi5462m&r57m;
wire cdxi8460m = cdxi5780m&r58m;
wire cdxi8461m = cdxi5424m&r59m;
wire cdxi8462m = cdxi5387m&r60m;
wire cdxi8463m = cdxi5349m&r61m;
wire cdxi8464m = cdxi5311m&r62m;
wire cdxi8465m = cdxi5154m&r83m;
wire cdxi8466m = cdxi4991m&r84m;
wire cdxi8467m = cdxi5136m&r85m;
wire cdxi8468m = cdxi5064m&r86m;
wire cdxi8469m = cdxi4973m&r87m;
wire cdxi8470m = cdxi4953m&r88m;
wire cdxi8471m = cdxi4934m&r89m;
wire cdxi8472m = cdxi5101m&r90m;
wire cdxi8473m = cdxi5083m&r91m;
wire cdxi8474m = cdxi4915m&r92m;
wire cdxi8475m = cdxi5065m&r93m;
wire cdxi8476m = cdxi4895m&r94m;
wire cdxi8477m = cdxi5028m&r95m;
wire cdxi8478m = cdxi5009m&r96m;
wire cdxi8479m = cdxi4873m&r97m;
wire cdxi8480m = cdxi4732m&r113m;
wire cdxi8481m = cdxi4742m&r114m;
wire cdxi8482m = cdxi4762m&r115m;
wire cdxi8483m = cdxi4722m&r116m;
wire cdxi8484m = cdxi4711m&r117m;
wire cdxi8485m = cdxi4743m&r118m;
wire cdxi8486m = (cdxi125m ^ cdxi8424m ^ cdxi8425m ^ cdxi8426m ^ cdxi8427m ^ cdxi8428m ^ cdxi8429m ^ cdxi8430m ^ cdxi8431m ^ cdxi8432m ^ cdxi8433m ^ cdxi8434m ^ cdxi8435m ^ cdxi8436m ^ cdxi8437m ^ cdxi8438m ^ cdxi8439m ^ cdxi8440m ^ cdxi8441m ^ cdxi8442m ^ cdxi8443m ^ cdxi8444m ^ cdxi8445m ^ cdxi8446m ^ cdxi8447m ^ cdxi8448m ^ cdxi8449m ^ cdxi8450m ^ cdxi8451m ^ cdxi8452m ^ cdxi8453m ^ cdxi8454m ^ cdxi8455m ^ cdxi8456m ^ cdxi8457m ^ cdxi8458m ^ cdxi8459m ^ cdxi8460m ^ cdxi8461m ^ cdxi8462m ^ cdxi8463m ^ cdxi8464m ^ cdxi8465m ^ cdxi8466m ^ cdxi8467m ^ cdxi8468m ^ cdxi8469m ^ cdxi8470m ^ cdxi8471m ^ cdxi8472m ^ cdxi8473m ^ cdxi8474m ^ cdxi8475m ^ cdxi8476m ^ cdxi8477m ^ cdxi8478m ^ cdxi8479m ^ cdxi8480m ^ cdxi8481m ^ cdxi8482m ^ cdxi8483m ^ cdxi8484m ^ cdxi8485m);
wire cdxi8487m = a1&cdxi8486m;
wire cdxi8488m = (reg_1_133);
wire cdxi8489m = reg_1_3&cdxi7079m;
wire cdxi8490m = reg_1_2&cdxi7145m;
wire cdxi8491m = reg_1_2&cdxi7146m;
wire cdxi8492m = reg_1_2&cdxi7147m;
wire cdxi8493m = reg_1_2&cdxi7148m;
wire cdxi8494m = reg_1_2&cdxi7149m;
wire cdxi8495m = reg_1_4&cdxi7219m;
wire cdxi8496m = reg_1_3&cdxi7084m;
wire cdxi8497m = reg_1_3&cdxi7085m;
wire cdxi8498m = reg_1_3&cdxi7086m;
wire cdxi8499m = reg_1_3&cdxi7087m;
wire cdxi8500m = reg_1_2&cdxi7150m;
wire cdxi8501m = reg_1_2&cdxi7151m;
wire cdxi8502m = reg_1_2&cdxi7152m;
wire cdxi8503m = reg_1_2&cdxi7153m;
wire cdxi8504m = reg_1_2&cdxi7154m;
wire cdxi8505m = reg_1_2&cdxi7155m;
wire cdxi8506m = reg_1_2&cdxi7156m;
wire cdxi8507m = reg_1_2&cdxi7157m;
wire cdxi8508m = reg_1_2&cdxi7158m;
wire cdxi8509m = reg_1_2&cdxi7159m;
wire cdxi8510m = reg_1_5&cdxi7029m;
wire cdxi8511m = reg_1_4&cdxi7229m;
wire cdxi8512m = reg_1_4&cdxi7230m;
wire cdxi8513m = reg_1_4&cdxi7231m;
wire cdxi8514m = reg_1_3&cdxi7094m;
wire cdxi8515m = reg_1_3&cdxi7095m;
wire cdxi8516m = reg_1_3&cdxi7096m;
wire cdxi8517m = reg_1_3&cdxi7097m;
wire cdxi8518m = reg_1_3&cdxi7098m;
wire cdxi8519m = reg_1_3&cdxi7099m;
wire cdxi8520m = reg_1_2&cdxi7160m;
wire cdxi8521m = reg_1_2&cdxi7161m;
wire cdxi8522m = reg_1_2&cdxi7162m;
wire cdxi8523m = reg_1_2&cdxi7163m;
wire cdxi8524m = reg_1_2&cdxi7164m;
wire cdxi8525m = reg_1_2&cdxi7165m;
wire cdxi8526m = reg_1_2&cdxi7166m;
wire cdxi8527m = reg_1_2&cdxi7167m;
wire cdxi8528m = reg_1_2&cdxi7168m;
wire cdxi8529m = reg_1_2&cdxi7169m;
wire cdxi8530m = reg_1_6&cdxi6972m;
wire cdxi8531m = reg_1_5&cdxi7039m;
wire cdxi8532m = reg_1_5&cdxi7040m;
wire cdxi8533m = reg_1_4&cdxi7239m;
wire cdxi8534m = reg_1_4&cdxi7240m;
wire cdxi8535m = reg_1_4&cdxi7241m;
wire cdxi8536m = reg_1_3&cdxi7104m;
wire cdxi8537m = reg_1_3&cdxi7105m;
wire cdxi8538m = reg_1_3&cdxi7106m;
wire cdxi8539m = reg_1_3&cdxi7107m;
wire cdxi8540m = reg_1_2&cdxi7170m;
wire cdxi8541m = reg_1_2&cdxi7171m;
wire cdxi8542m = reg_1_2&cdxi7172m;
wire cdxi8543m = reg_1_2&cdxi7173m;
wire cdxi8544m = reg_1_2&cdxi7174m;
wire cdxi8545m = reg_1_7&cdxi8259m;
wire cdxi8546m = reg_1_6&cdxi6946m;
wire cdxi8547m = reg_1_5&cdxi7013m;
wire cdxi8548m = reg_1_4&cdxi7213m;
wire cdxi8549m = reg_1_3&cdxi7078m;
wire cdxi8550m = reg_1_2&cdxi7144m;
wire cdxi8551m = (cdxi8489m ^ cdxi8490m ^ cdxi8491m ^ cdxi8492m ^ cdxi8493m ^ cdxi8494m ^ cdxi8495m ^ cdxi8496m ^ cdxi8497m ^ cdxi8498m ^ cdxi8499m ^ cdxi8500m ^ cdxi8501m ^ cdxi8502m ^ cdxi8503m ^ cdxi8504m ^ cdxi8505m ^ cdxi8506m ^ cdxi8507m ^ cdxi8508m ^ cdxi8509m ^ cdxi8510m ^ cdxi8511m ^ cdxi8512m ^ cdxi8513m ^ cdxi8514m ^ cdxi8515m ^ cdxi8516m ^ cdxi8517m ^ cdxi8518m ^ cdxi8519m ^ cdxi8520m ^ cdxi8521m ^ cdxi8522m ^ cdxi8523m ^ cdxi8524m ^ cdxi8525m ^ cdxi8526m ^ cdxi8527m ^ cdxi8528m ^ cdxi8529m ^ cdxi8530m ^ cdxi8531m ^ cdxi8532m ^ cdxi8533m ^ cdxi8534m ^ cdxi8535m ^ cdxi8536m ^ cdxi8537m ^ cdxi8538m ^ cdxi8539m ^ cdxi8540m ^ cdxi8541m ^ cdxi8542m ^ cdxi8543m ^ cdxi8544m ^ cdxi8545m ^ cdxi8546m ^ cdxi8547m ^ cdxi8548m ^ cdxi8549m ^ cdxi8550m ^ cdxi8488m);
wire cdxi8552m = reg_1_0&cdxi8551m;
wire cdxi8553m = cdxi4712m ^ cdxi4711m ^ cdxi4762m ^ cdxi4742m;
wire cdxi8554m = cdxi4712m&cdxi4m;
wire cdxi8555m = reg_1_1&cdxi4685m;
wire cdxi8556m = cdxi4743m&cdxi6m;
wire cdxi8557m = reg_1_2&cdxi4699m;
wire cdxi8558m = cdxi4711m&cdxi6m;
wire cdxi8559m = reg_1_3&cdxi4699m;
wire cdxi8560m = cdxi4711m&r1m;
wire cdxi8561m = cdxi4743m&r2m;
wire cdxi8562m = (cdxi13m ^ cdxi8560m ^ cdxi8561m);
wire cdxi8563m = cdxi4712m&cdxi8562m;
wire cdxi8564m = reg_1_3&cdxi4669m;
wire cdxi8565m = reg_1_2&cdxi4674m;
wire cdxi8566m = (cdxi8564m ^ cdxi8565m ^ cdxi4885m);
wire cdxi8567m = reg_1_1&cdxi8566m;
wire cdxi8568m = cdxi4712m&cdxi4746m;
wire cdxi8569m = reg_1_1&cdxi4751m;
wire cdxi8570m = cdxi4712m&cdxi4828m;
wire cdxi8571m = reg_1_1&cdxi4833m;
wire cdxi8572m = cdxi4712m&cdxi4783m;
wire cdxi8573m = reg_1_1&cdxi4788m;
wire cdxi8574m = cdxi4712m&cdxi4852m;
wire cdxi8575m = reg_1_1&cdxi4857m;
wire cdxi8576m = cdxi4722m&cdxi4852m;
wire cdxi8577m = reg_1_4&cdxi4857m;
wire cdxi8578m = cdxi5136m&r0m;
wire cdxi8579m = cdxi4712m&cdxi4772m;
wire cdxi8580m = cdxi4712m&cdxi4773m;
wire cdxi8581m = cdxi4742m&r10m;
wire cdxi8582m = cdxi4762m&r11m;
wire cdxi8583m = cdxi4712m&r25m;
wire cdxi8584m = (cdxi40m ^ cdxi8578m ^ cdxi8579m ^ cdxi8580m ^ cdxi8581m ^ cdxi8582m ^ cdxi8583m);
wire cdxi8585m = a1&cdxi8584m;
wire cdxi8586m = reg_1_5&reg_1_6&cdxi4664m;
wire cdxi8587m = reg_1_1&cdxi4777m;
wire cdxi8588m = reg_1_1&cdxi4778m;
wire cdxi8589m = reg_1_6&cdxi4963m;
wire cdxi8590m = reg_1_5&cdxi4905m;
wire cdxi8591m = reg_1_1&cdxi4776m;
wire cdxi8592m = (cdxi8586m ^ cdxi8587m ^ cdxi8588m ^ cdxi8589m ^ cdxi8590m ^ cdxi8591m ^ cdxi5515m);
wire cdxi8593m = reg_1_0&cdxi8592m;
wire cdxi8594m = cdxi4742m&cdxi4733m;
wire cdxi8595m = cdxi4712m&cdxi4850m;
wire cdxi8596m = cdxi4712m&cdxi4851m;
wire cdxi8597m = cdxi4732m&r11m;
wire cdxi8598m = cdxi4742m&r12m;
wire cdxi8599m = cdxi4712m&r27m;
wire cdxi8600m = (cdxi42m ^ cdxi8594m ^ cdxi8595m ^ cdxi8596m ^ cdxi8597m ^ cdxi8598m ^ cdxi8599m);
wire cdxi8601m = a1&cdxi8600m;
wire cdxi8602m = reg_1_6&cdxi4738m;
wire cdxi8603m = reg_1_1&cdxi4855m;
wire cdxi8604m = reg_1_1&cdxi4856m;
wire cdxi8605m = reg_1_7&cdxi4905m;
wire cdxi8606m = reg_1_6&cdxi4737m;
wire cdxi8607m = reg_1_1&cdxi4854m;
wire cdxi8608m = (cdxi8602m ^ cdxi8603m ^ cdxi8604m ^ cdxi8605m ^ cdxi8606m ^ cdxi8607m ^ cdxi5551m);
wire cdxi8609m = reg_1_0&cdxi8608m;
wire cdxi8610m = a1&cdxi5178m;
wire cdxi8611m = reg_1_0&cdxi5187m;
wire cdxi8612m = a1&cdxi5216m;
wire cdxi8613m = reg_1_0&cdxi5225m;
wire cdxi8614m = cdxi4712m&cdxi8001m;
wire cdxi8615m = reg_1_1&cdxi8009m;
wire cdxi8616m = cdxi4712m&cdxi5298m;
wire cdxi8617m = reg_1_1&cdxi5307m;
wire cdxi8618m = cdxi5950m&r0m;
wire cdxi8619m = cdxi4954m&cdxi4817m;
wire cdxi8620m = cdxi4916m&cdxi4772m;
wire cdxi8621m = cdxi4916m&cdxi4773m;
wire cdxi8622m = cdxi4762m&cdxi4977m;
wire cdxi8623m = cdxi4973m&r10m;
wire cdxi8624m = cdxi4953m&r11m;
wire cdxi8625m = cdxi4896m&r22m;
wire cdxi8626m = cdxi4954m&r23m;
wire cdxi8627m = cdxi4916m&r25m;
wire cdxi8628m = cdxi4742m&r37m;
wire cdxi8629m = cdxi4762m&r38m;
wire cdxi8630m = cdxi4722m&r40m;
wire cdxi8631m = cdxi4712m&r59m;
wire cdxi8632m = (cdxi79m ^ cdxi8618m ^ cdxi8619m ^ cdxi8620m ^ cdxi8621m ^ cdxi8622m ^ cdxi8623m ^ cdxi8624m ^ cdxi8625m ^ cdxi8626m ^ cdxi8627m ^ cdxi8628m ^ cdxi8629m ^ cdxi8630m ^ cdxi8631m);
wire cdxi8633m = a1&cdxi8632m;
wire cdxi8634m = reg_1_4&cdxi8586m;
wire cdxi8635m = reg_1_1&cdxi5146m;
wire cdxi8636m = reg_1_1&cdxi5147m;
wire cdxi8637m = reg_1_1&cdxi5148m;
wire cdxi8638m = reg_1_5&cdxi4986m;
wire cdxi8639m = reg_1_4&cdxi8589m;
wire cdxi8640m = reg_1_4&cdxi8590m;
wire cdxi8641m = reg_1_1&cdxi5149m;
wire cdxi8642m = reg_1_1&cdxi5150m;
wire cdxi8643m = reg_1_1&cdxi5151m;
wire cdxi8644m = reg_1_6&cdxi4964m;
wire cdxi8645m = reg_1_5&cdxi4982m;
wire cdxi8646m = reg_1_4&cdxi5515m;
wire cdxi8647m = reg_1_1&cdxi5145m;
wire cdxi8648m = (cdxi8634m ^ cdxi8635m ^ cdxi8636m ^ cdxi8637m ^ cdxi8638m ^ cdxi8639m ^ cdxi8640m ^ cdxi8641m ^ cdxi8642m ^ cdxi8643m ^ cdxi8644m ^ cdxi8645m ^ cdxi8646m ^ cdxi8647m ^ cdxi6538m);
wire cdxi8649m = reg_1_0&cdxi8648m;
wire cdxi8650m = a1&cdxi6100m;
wire cdxi8651m = reg_1_0&cdxi6117m;
wire cdxi8652m = cdxi4712m&cdxi5965m;
wire cdxi8653m = reg_1_1&cdxi5982m;
wire cdxi8654m = cdxi4712m&cdxi8095m;
wire cdxi8655m = reg_1_1&cdxi8111m;
wire cdxi8656m = cdxi4712m&cdxi6166m;
wire cdxi8657m = reg_1_1&cdxi6183m;
wire cdxi8658m = cdxi5848m&cdxi4733m;
wire cdxi8659m = cdxi5498m&cdxi4753m;
wire cdxi8660m = cdxi4874m&cdxi5155m;
wire cdxi8661m = cdxi4874m&cdxi5156m;
wire cdxi8662m = cdxi4874m&cdxi5157m;
wire cdxi8663m = cdxi5136m&cdxi4939m;
wire cdxi8664m = cdxi5101m&cdxi4995m;
wire cdxi8665m = cdxi5640m&r11m;
wire cdxi8666m = cdxi5848m&r12m;
wire cdxi8667m = cdxi4896m&cdxi5122m;
wire cdxi8668m = cdxi5641m&r20m;
wire cdxi8669m = cdxi5498m&r21m;
wire cdxi8670m = cdxi4874m&cdxi5158m;
wire cdxi8671m = cdxi4874m&cdxi5159m;
wire cdxi8672m = cdxi4874m&cdxi5160m;
wire cdxi8673m = cdxi5154m&r34m;
wire cdxi8674m = cdxi4991m&r35m;
wire cdxi8675m = cdxi5136m&r36m;
wire cdxi8676m = cdxi4934m&r40m;
wire cdxi8677m = cdxi5101m&r41m;
wire cdxi8678m = cdxi5083m&r42m;
wire cdxi8679m = cdxi4935m&r56m;
wire cdxi8680m = cdxi4896m&r57m;
wire cdxi8681m = cdxi4954m&r58m;
wire cdxi8682m = cdxi4874m&r62m;
wire cdxi8683m = cdxi4732m&r76m;
wire cdxi8684m = cdxi4742m&r77m;
wire cdxi8685m = cdxi4762m&r78m;
wire cdxi8686m = cdxi4711m&r82m;
wire cdxi8687m = cdxi4712m&r96m;
wire cdxi8688m = (cdxi111m ^ cdxi8658m ^ cdxi8659m ^ cdxi8660m ^ cdxi8661m ^ cdxi8662m ^ cdxi8663m ^ cdxi8664m ^ cdxi8665m ^ cdxi8666m ^ cdxi8667m ^ cdxi8668m ^ cdxi8669m ^ cdxi8670m ^ cdxi8671m ^ cdxi8672m ^ cdxi8673m ^ cdxi8674m ^ cdxi8675m ^ cdxi8676m ^ cdxi8677m ^ cdxi8678m ^ cdxi8679m ^ cdxi8680m ^ cdxi8681m ^ cdxi8682m ^ cdxi8683m ^ cdxi8684m ^ cdxi8685m ^ cdxi8686m ^ cdxi8687m);
wire cdxi8689m = a1&cdxi8688m;
wire cdxi8690m = reg_1_3&cdxi8065m;
wire cdxi8691m = reg_1_1&cdxi6035m;
wire cdxi8692m = reg_1_1&cdxi6036m;
wire cdxi8693m = reg_1_1&cdxi6037m;
wire cdxi8694m = reg_1_1&cdxi6038m;
wire cdxi8695m = reg_1_5&cdxi5698m;
wire cdxi8696m = reg_1_3&cdxi8069m;
wire cdxi8697m = reg_1_3&cdxi8070m;
wire cdxi8698m = reg_1_3&cdxi8071m;
wire cdxi8699m = reg_1_1&cdxi6039m;
wire cdxi8700m = reg_1_1&cdxi6040m;
wire cdxi8701m = reg_1_1&cdxi6041m;
wire cdxi8702m = reg_1_1&cdxi6042m;
wire cdxi8703m = reg_1_1&cdxi6043m;
wire cdxi8704m = reg_1_1&cdxi6044m;
wire cdxi8705m = reg_1_6&cdxi5669m;
wire cdxi8706m = reg_1_5&cdxi5704m;
wire cdxi8707m = reg_1_5&cdxi5705m;
wire cdxi8708m = reg_1_3&cdxi8075m;
wire cdxi8709m = reg_1_3&cdxi8076m;
wire cdxi8710m = reg_1_3&cdxi8077m;
wire cdxi8711m = reg_1_1&cdxi6045m;
wire cdxi8712m = reg_1_1&cdxi6046m;
wire cdxi8713m = reg_1_1&cdxi6047m;
wire cdxi8714m = reg_1_1&cdxi6048m;
wire cdxi8715m = reg_1_7&cdxi6400m;
wire cdxi8716m = reg_1_6&cdxi5658m;
wire cdxi8717m = reg_1_5&cdxi5693m;
wire cdxi8718m = reg_1_3&cdxi6677m;
wire cdxi8719m = reg_1_1&cdxi6034m;
wire cdxi8720m = (cdxi8690m ^ cdxi8691m ^ cdxi8692m ^ cdxi8693m ^ cdxi8694m ^ cdxi8695m ^ cdxi8696m ^ cdxi8697m ^ cdxi8698m ^ cdxi8699m ^ cdxi8700m ^ cdxi8701m ^ cdxi8702m ^ cdxi8703m ^ cdxi8704m ^ cdxi8705m ^ cdxi8706m ^ cdxi8707m ^ cdxi8708m ^ cdxi8709m ^ cdxi8710m ^ cdxi8711m ^ cdxi8712m ^ cdxi8713m ^ cdxi8714m ^ cdxi8715m ^ cdxi8716m ^ cdxi8717m ^ cdxi8718m ^ cdxi8719m ^ cdxi7456m);
wire cdxi8721m = reg_1_0&cdxi8720m;
wire cdxi8722m = cdxi4712m&cdxi7076m;
wire cdxi8723m = reg_1_1&cdxi7109m;
wire cdxi8724m = cdxi4743m&cdxi7142m;
wire cdxi8725m = reg_1_2&cdxi7175m;
wire cdxi8726m = cdxi4873m&cdxi5712m;
wire cdxi8727m = cdxi4874m&cdxi5984m;
wire cdxi8728m = cdxi4875m&cdxi6086m;
wire cdxi8729m = cdxi5314m&cdxi5292m;
wire cdxi8730m = cdxi5314m&cdxi5293m;
wire cdxi8731m = cdxi5314m&cdxi5294m;
wire cdxi8732m = cdxi6778m&r7m;
wire cdxi8733m = cdxi5780m&cdxi4939m;
wire cdxi8734m = cdxi4873m&cdxi5716m;
wire cdxi8735m = cdxi5311m&cdxi4995m;
wire cdxi8736m = cdxi4873m&cdxi5718m;
wire cdxi8737m = cdxi4916m&cdxi5888m;
wire cdxi8738m = cdxi4874m&cdxi5988m;
wire cdxi8739m = cdxi4874m&cdxi5989m;
wire cdxi8740m = cdxi4874m&cdxi5990m;
wire cdxi8741m = cdxi4875m&cdxi6090m;
wire cdxi8742m = cdxi4875m&cdxi6091m;
wire cdxi8743m = cdxi4875m&cdxi6092m;
wire cdxi8744m = cdxi5314m&cdxi5295m;
wire cdxi8745m = cdxi5314m&cdxi5296m;
wire cdxi8746m = cdxi5314m&cdxi5297m;
wire cdxi8747m = cdxi4953m&cdxi5437m;
wire cdxi8748m = cdxi5640m&r29m;
wire cdxi8749m = cdxi5604m&r30m;
wire cdxi8750m = cdxi5779m&r32m;
wire cdxi8751m = cdxi5883m&r33m;
wire cdxi8752m = cdxi5009m&cdxi5652m;
wire cdxi8753m = cdxi5780m&r36m;
wire cdxi8754m = cdxi5424m&r37m;
wire cdxi8755m = cdxi5349m&r39m;
wire cdxi8756m = cdxi5311m&r41m;
wire cdxi8757m = cdxi5641m&r43m;
wire cdxi8758m = cdxi5605m&r44m;
wire cdxi8759m = cdxi5711m&r46m;
wire cdxi8760m = cdxi5425m&r47m;
wire cdxi8761m = cdxi5350m&r49m;
wire cdxi8762m = cdxi5312m&r51m;
wire cdxi8763m = cdxi5426m&r53m;
wire cdxi8764m = cdxi5351m&r55m;
wire cdxi8765m = cdxi5313m&r57m;
wire cdxi8766m = cdxi5314m&r60m;
wire cdxi8767m = cdxi4991m&r63m;
wire cdxi8768m = cdxi5064m&r64m;
wire cdxi8769m = cdxi4953m&r66m;
wire cdxi8770m = cdxi4934m&r67m;
wire cdxi8771m = cdxi5083m&r69m;
wire cdxi8772m = cdxi4915m&r71m;
wire cdxi8773m = cdxi5065m&r73m;
wire cdxi8774m = cdxi5028m&r75m;
wire cdxi8775m = cdxi5009m&r77m;
wire cdxi8776m = cdxi4873m&r80m;
wire cdxi8777m = cdxi4935m&r83m;
wire cdxi8778m = cdxi4954m&r85m;
wire cdxi8779m = cdxi4916m&r87m;
wire cdxi8780m = cdxi4874m&r90m;
wire cdxi8781m = cdxi4875m&r94m;
wire cdxi8782m = cdxi4732m&r98m;
wire cdxi8783m = cdxi4762m&r100m;
wire cdxi8784m = cdxi4722m&r102m;
wire cdxi8785m = cdxi4711m&r105m;
wire cdxi8786m = cdxi4743m&r109m;
wire cdxi8787m = cdxi4712m&r114m;
wire cdxi8788m = (cdxi120m ^ cdxi8726m ^ cdxi8727m ^ cdxi8728m ^ cdxi8729m ^ cdxi8730m ^ cdxi8731m ^ cdxi8732m ^ cdxi8733m ^ cdxi8734m ^ cdxi8735m ^ cdxi8736m ^ cdxi8737m ^ cdxi8738m ^ cdxi8739m ^ cdxi8740m ^ cdxi8741m ^ cdxi8742m ^ cdxi8743m ^ cdxi8744m ^ cdxi8745m ^ cdxi8746m ^ cdxi8747m ^ cdxi8748m ^ cdxi8749m ^ cdxi8750m ^ cdxi8751m ^ cdxi8752m ^ cdxi8753m ^ cdxi8754m ^ cdxi8755m ^ cdxi8756m ^ cdxi8757m ^ cdxi8758m ^ cdxi8759m ^ cdxi8760m ^ cdxi8761m ^ cdxi8762m ^ cdxi8763m ^ cdxi8764m ^ cdxi8765m ^ cdxi8766m ^ cdxi8767m ^ cdxi8768m ^ cdxi8769m ^ cdxi8770m ^ cdxi8771m ^ cdxi8772m ^ cdxi8773m ^ cdxi8774m ^ cdxi8775m ^ cdxi8776m ^ cdxi8777m ^ cdxi8778m ^ cdxi8779m ^ cdxi8780m ^ cdxi8781m ^ cdxi8782m ^ cdxi8783m ^ cdxi8784m ^ cdxi8785m ^ cdxi8786m ^ cdxi8787m);
wire cdxi8789m = a1&cdxi8788m;
wire cdxi8790m = (reg_1_128);
wire cdxi8791m = reg_1_2&cdxi6814m;
wire cdxi8792m = reg_1_1&cdxi6947m;
wire cdxi8793m = reg_1_1&cdxi6948m;
wire cdxi8794m = reg_1_1&cdxi6949m;
wire cdxi8795m = reg_1_1&cdxi6950m;
wire cdxi8796m = reg_1_1&cdxi6951m;
wire cdxi8797m = reg_1_3&reg_1_4&reg_1_5&cdxi7890m;
wire cdxi8798m = reg_1_2&cdxi6819m;
wire cdxi8799m = reg_1_2&cdxi6820m;
wire cdxi8800m = reg_1_2&cdxi6821m;
wire cdxi8801m = reg_1_2&cdxi6822m;
wire cdxi8802m = reg_1_1&cdxi6952m;
wire cdxi8803m = reg_1_1&cdxi6953m;
wire cdxi8804m = reg_1_1&cdxi6954m;
wire cdxi8805m = reg_1_1&cdxi6955m;
wire cdxi8806m = reg_1_1&cdxi6956m;
wire cdxi8807m = reg_1_1&cdxi6957m;
wire cdxi8808m = reg_1_1&cdxi6958m;
wire cdxi8809m = reg_1_1&cdxi6959m;
wire cdxi8810m = reg_1_1&cdxi6960m;
wire cdxi8811m = reg_1_1&cdxi6961m;
wire cdxi8812m = reg_1_4&cdxi6487m;
wire cdxi8813m = reg_1_3&reg_1_5&cdxi8043m;
wire cdxi8814m = reg_1_3&reg_1_4&reg_1_7&cdxi5368m;
wire cdxi8815m = reg_1_3&reg_1_4&reg_1_5&cdxi5443m;
wire cdxi8816m = reg_1_2&cdxi6829m;
wire cdxi8817m = reg_1_2&cdxi6830m;
wire cdxi8818m = reg_1_2&cdxi6831m;
wire cdxi8819m = reg_1_2&cdxi6832m;
wire cdxi8820m = reg_1_2&cdxi6833m;
wire cdxi8821m = reg_1_2&cdxi6834m;
wire cdxi8822m = reg_1_1&cdxi6962m;
wire cdxi8823m = reg_1_1&cdxi6963m;
wire cdxi8824m = reg_1_1&cdxi6964m;
wire cdxi8825m = reg_1_1&cdxi6965m;
wire cdxi8826m = reg_1_1&cdxi6966m;
wire cdxi8827m = reg_1_1&cdxi6967m;
wire cdxi8828m = reg_1_1&cdxi6968m;
wire cdxi8829m = reg_1_1&cdxi6969m;
wire cdxi8830m = reg_1_1&cdxi6970m;
wire cdxi8831m = reg_1_1&cdxi6971m;
wire cdxi8832m = reg_1_5&reg_1_7&cdxi5332m;
wire cdxi8833m = reg_1_4&cdxi6497m;
wire cdxi8834m = reg_1_4&cdxi6498m;
wire cdxi8835m = reg_1_3&reg_1_7&cdxi6261m;
wire cdxi8836m = reg_1_3&reg_1_5&cdxi6608m;
wire cdxi8837m = reg_1_3&reg_1_4&cdxi6470m;
wire cdxi8838m = reg_1_2&cdxi6839m;
wire cdxi8839m = reg_1_2&cdxi6840m;
wire cdxi8840m = reg_1_2&cdxi6841m;
wire cdxi8841m = reg_1_2&cdxi6842m;
wire cdxi8842m = reg_1_1&cdxi6972m;
wire cdxi8843m = reg_1_1&cdxi6973m;
wire cdxi8844m = reg_1_1&cdxi6974m;
wire cdxi8845m = reg_1_1&cdxi6975m;
wire cdxi8846m = reg_1_1&cdxi6976m;
wire cdxi8847m = reg_1_7&cdxi6263m;
wire cdxi8848m = reg_1_5&cdxi7319m;
wire cdxi8849m = reg_1_4&cdxi6471m;
wire cdxi8850m = reg_1_3&cdxi7590m;
wire cdxi8851m = reg_1_2&cdxi6813m;
wire cdxi8852m = reg_1_1&cdxi6946m;
wire cdxi8853m = (cdxi8791m ^ cdxi8792m ^ cdxi8793m ^ cdxi8794m ^ cdxi8795m ^ cdxi8796m ^ cdxi8797m ^ cdxi8798m ^ cdxi8799m ^ cdxi8800m ^ cdxi8801m ^ cdxi8802m ^ cdxi8803m ^ cdxi8804m ^ cdxi8805m ^ cdxi8806m ^ cdxi8807m ^ cdxi8808m ^ cdxi8809m ^ cdxi8810m ^ cdxi8811m ^ cdxi8812m ^ cdxi8813m ^ cdxi8814m ^ cdxi8815m ^ cdxi8816m ^ cdxi8817m ^ cdxi8818m ^ cdxi8819m ^ cdxi8820m ^ cdxi8821m ^ cdxi8822m ^ cdxi8823m ^ cdxi8824m ^ cdxi8825m ^ cdxi8826m ^ cdxi8827m ^ cdxi8828m ^ cdxi8829m ^ cdxi8830m ^ cdxi8831m ^ cdxi8832m ^ cdxi8833m ^ cdxi8834m ^ cdxi8835m ^ cdxi8836m ^ cdxi8837m ^ cdxi8838m ^ cdxi8839m ^ cdxi8840m ^ cdxi8841m ^ cdxi8842m ^ cdxi8843m ^ cdxi8844m ^ cdxi8845m ^ cdxi8846m ^ cdxi8847m ^ cdxi8848m ^ cdxi8849m ^ cdxi8850m ^ cdxi8851m ^ cdxi8852m ^ cdxi8790m);
wire cdxi8854m = reg_1_0&cdxi8853m;
wire cdxi8855m = cdxi4712m&cdxi8486m;
wire cdxi8856m = reg_1_1&cdxi8551m;
wire cdxi8857m = 0&0 ^ cdxi4712m ^ cdxi4722m ^ cdxi4742m ^ cdxi4732m;
wire cdxi8858m = cdxi4712m&cdxi4755m;
wire cdxi8859m = reg_1_1&cdxi4760m;
wire cdxi8860m = cdxi4712m&cdxi4765m;
wire cdxi8861m = reg_1_1&cdxi4770m;
wire cdxi8862m = cdxi4711m&cdxi4852m;
wire cdxi8863m = reg_1_3&cdxi4857m;
wire cdxi8864m = cdxi5028m&r0m;
wire cdxi8865m = cdxi4954m&r1m;
wire cdxi8866m = cdxi4875m&r4m;
wire cdxi8867m = cdxi4762m&r7m;
wire cdxi8868m = cdxi4743m&r10m;
wire cdxi8869m = cdxi4712m&r15m;
wire cdxi8870m = (cdxi30m ^ cdxi8864m ^ cdxi8865m ^ cdxi8866m ^ cdxi8867m ^ cdxi8868m ^ cdxi8869m);
wire cdxi8871m = a1&cdxi8870m;
wire cdxi8872m = reg_1_2&cdxi7815m;
wire cdxi8873m = reg_1_1&cdxi7831m;
wire cdxi8874m = reg_1_1&cdxi7832m;
wire cdxi8875m = reg_1_5&cdxi4884m;
wire cdxi8876m = reg_1_2&cdxi4963m;
wire cdxi8877m = reg_1_1&cdxi5037m;
wire cdxi8878m = (cdxi8872m ^ cdxi8873m ^ cdxi8874m ^ cdxi8875m ^ cdxi8876m ^ cdxi8877m ^ cdxi5368m);
wire cdxi8879m = reg_1_0&cdxi8878m;
wire cdxi8880m = cdxi4743m&cdxi4992m;
wire cdxi8881m = cdxi4954m&cdxi4790m;
wire cdxi8882m = cdxi4875m&cdxi4781m;
wire cdxi8883m = cdxi4875m&cdxi4782m;
wire cdxi8884m = cdxi4991m&r7m;
wire cdxi8885m = cdxi4743m&cdxi4995m;
wire cdxi8886m = cdxi4743m&cdxi4996m;
wire cdxi8887m = cdxi4935m&r15m;
wire cdxi8888m = cdxi4954m&r17m;
wire cdxi8889m = cdxi4875m&r26m;
wire cdxi8890m = cdxi4732m&r30m;
wire cdxi8891m = cdxi4762m&r32m;
wire cdxi8892m = cdxi4743m&r41m;
wire cdxi8893m = cdxi4712m&r51m;
wire cdxi8894m = (cdxi71m ^ cdxi8880m ^ cdxi8881m ^ cdxi8882m ^ cdxi8883m ^ cdxi8884m ^ cdxi8885m ^ cdxi8886m ^ cdxi8887m ^ cdxi8888m ^ cdxi8889m ^ cdxi8890m ^ cdxi8891m ^ cdxi8892m ^ cdxi8893m);
wire cdxi8895m = a1&cdxi8894m;
wire cdxi8896m = reg_1_2&cdxi5001m;
wire cdxi8897m = reg_1_1&cdxi5236m;
wire cdxi8898m = reg_1_1&cdxi5237m;
wire cdxi8899m = reg_1_1&cdxi5238m;
wire cdxi8900m = reg_1_5&cdxi7890m;
wire cdxi8901m = reg_1_2&cdxi5004m;
wire cdxi8902m = reg_1_2&cdxi5005m;
wire cdxi8903m = reg_1_1&cdxi5239m;
wire cdxi8904m = reg_1_1&cdxi5240m;
wire cdxi8905m = reg_1_1&cdxi5241m;
wire cdxi8906m = reg_1_7&cdxi5368m;
wire cdxi8907m = reg_1_5&cdxi5443m;
wire cdxi8908m = reg_1_2&cdxi5000m;
wire cdxi8909m = reg_1_1&cdxi5235m;
wire cdxi8910m = (cdxi8896m ^ cdxi8897m ^ cdxi8898m ^ cdxi8899m ^ cdxi8900m ^ cdxi8901m ^ cdxi8902m ^ cdxi8903m ^ cdxi8904m ^ cdxi8905m ^ cdxi8906m ^ cdxi8907m ^ cdxi8908m ^ cdxi8909m ^ cdxi6470m);
wire cdxi8911m = reg_1_0&cdxi8910m;
wire cdxi8912m = cdxi5779m&r0m;
wire cdxi8913m = cdxi4916m&cdxi4826m;
wire cdxi8914m = cdxi4874m&cdxi4763m;
wire cdxi8915m = cdxi4874m&cdxi4764m;
wire cdxi8916m = cdxi4953m&r8m;
wire cdxi8917m = cdxi4711m&cdxi4958m;
wire cdxi8918m = cdxi4915m&r10m;
wire cdxi8919m = cdxi4954m&r18m;
wire cdxi8920m = cdxi4916m&r19m;
wire cdxi8921m = cdxi4874m&r22m;
wire cdxi8922m = cdxi4762m&r33m;
wire cdxi8923m = cdxi4722m&r34m;
wire cdxi8924m = cdxi4711m&r37m;
wire cdxi8925m = cdxi4712m&r53m;
wire cdxi8926m = (cdxi73m ^ cdxi8912m ^ cdxi8913m ^ cdxi8914m ^ cdxi8915m ^ cdxi8916m ^ cdxi8917m ^ cdxi8918m ^ cdxi8919m ^ cdxi8920m ^ cdxi8921m ^ cdxi8922m ^ cdxi8923m ^ cdxi8924m ^ cdxi8925m);
wire cdxi8927m = a1&cdxi8926m;
wire cdxi8928m = reg_1_3&cdxi4965m;
wire cdxi8929m = reg_1_1&cdxi5093m;
wire cdxi8930m = reg_1_1&cdxi5094m;
wire cdxi8931m = reg_1_1&cdxi5095m;
wire cdxi8932m = reg_1_4&cdxi7906m;
wire cdxi8933m = reg_1_3&cdxi4968m;
wire cdxi8934m = reg_1_3&cdxi4969m;
wire cdxi8935m = reg_1_1&cdxi5096m;
wire cdxi8936m = reg_1_1&cdxi5097m;
wire cdxi8937m = reg_1_1&cdxi5098m;
wire cdxi8938m = reg_1_5&cdxi4925m;
wire cdxi8939m = reg_1_4&cdxi5369m;
wire cdxi8940m = reg_1_3&cdxi4964m;
wire cdxi8941m = reg_1_1&cdxi5092m;
wire cdxi8942m = (cdxi8928m ^ cdxi8929m ^ cdxi8930m ^ cdxi8931m ^ cdxi8932m ^ cdxi8933m ^ cdxi8934m ^ cdxi8935m ^ cdxi8936m ^ cdxi8937m ^ cdxi8938m ^ cdxi8939m ^ cdxi8940m ^ cdxi8941m ^ cdxi6262m);
wire cdxi8943m = reg_1_0&cdxi8942m;
wire cdxi8944m = a1&cdxi6065m;
wire cdxi8945m = reg_1_0&cdxi6082m;
wire cdxi8946m = a1&cdxi6166m;
wire cdxi8947m = reg_1_0&cdxi6183m;
wire cdxi8948m = cdxi5311m&cdxi4733m;
wire cdxi8949m = cdxi4874m&cdxi5066m;
wire cdxi8950m = cdxi4875m&cdxi5269m;
wire cdxi8951m = cdxi5314m&cdxi4839m;
wire cdxi8952m = cdxi5314m&cdxi4840m;
wire cdxi8953m = cdxi5604m&r7m;
wire cdxi8954m = cdxi5009m&cdxi4939m;
wire cdxi8955m = cdxi5424m&r9m;
wire cdxi8956m = cdxi5311m&r12m;
wire cdxi8957m = cdxi5605m&r13m;
wire cdxi8958m = cdxi4874m&cdxi5069m;
wire cdxi8959m = cdxi4874m&cdxi5070m;
wire cdxi8960m = cdxi4875m&cdxi5272m;
wire cdxi8961m = cdxi4875m&cdxi5273m;
wire cdxi8962m = cdxi5314m&r24m;
wire cdxi8963m = cdxi5064m&r28m;
wire cdxi8964m = cdxi4934m&r29m;
wire cdxi8965m = cdxi4915m&r32m;
wire cdxi8966m = cdxi5065m&r33m;
wire cdxi8967m = cdxi5009m&r36m;
wire cdxi8968m = cdxi4873m&r39m;
wire cdxi8969m = cdxi4935m&r43m;
wire cdxi8970m = cdxi4916m&r46m;
wire cdxi8971m = cdxi4874m&r49m;
wire cdxi8972m = cdxi4875m&r55m;
wire cdxi8973m = cdxi4732m&r63m;
wire cdxi8974m = cdxi4722m&r66m;
wire cdxi8975m = cdxi4711m&r69m;
wire cdxi8976m = cdxi4743m&r75m;
wire cdxi8977m = cdxi4712m&r85m;
wire cdxi8978m = (cdxi100m ^ cdxi8948m ^ cdxi8949m ^ cdxi8950m ^ cdxi8951m ^ cdxi8952m ^ cdxi8953m ^ cdxi8954m ^ cdxi8955m ^ cdxi8956m ^ cdxi8957m ^ cdxi8958m ^ cdxi8959m ^ cdxi8960m ^ cdxi8961m ^ cdxi8962m ^ cdxi8963m ^ cdxi8964m ^ cdxi8965m ^ cdxi8966m ^ cdxi8967m ^ cdxi8968m ^ cdxi8969m ^ cdxi8970m ^ cdxi8971m ^ cdxi8972m ^ cdxi8973m ^ cdxi8974m ^ cdxi8975m ^ cdxi8976m ^ cdxi8977m);
wire cdxi8979m = a1&cdxi8978m;
wire cdxi8980m = reg_1_2&cdxi5624m;
wire cdxi8981m = reg_1_1&cdxi5832m;
wire cdxi8982m = reg_1_1&cdxi5833m;
wire cdxi8983m = reg_1_1&cdxi5834m;
wire cdxi8984m = reg_1_1&cdxi5835m;
wire cdxi8985m = reg_1_3&cdxi8037m;
wire cdxi8986m = reg_1_2&cdxi5628m;
wire cdxi8987m = reg_1_2&cdxi5629m;
wire cdxi8988m = reg_1_2&cdxi5630m;
wire cdxi8989m = reg_1_1&cdxi5836m;
wire cdxi8990m = reg_1_1&cdxi5837m;
wire cdxi8991m = reg_1_1&cdxi5838m;
wire cdxi8992m = reg_1_1&cdxi5839m;
wire cdxi8993m = reg_1_1&cdxi5840m;
wire cdxi8994m = reg_1_1&cdxi5841m;
wire cdxi8995m = reg_1_4&cdxi5456m;
wire cdxi8996m = reg_1_3&cdxi8043m;
wire cdxi8997m = reg_1_3&cdxi8044m;
wire cdxi8998m = reg_1_2&cdxi5634m;
wire cdxi8999m = reg_1_2&cdxi5635m;
wire cdxi9000m = reg_1_2&cdxi5636m;
wire cdxi9001m = reg_1_1&cdxi5842m;
wire cdxi9002m = reg_1_1&cdxi5843m;
wire cdxi9003m = reg_1_1&cdxi5844m;
wire cdxi9004m = reg_1_1&cdxi5845m;
wire cdxi9005m = reg_1_7&cdxi5332m;
wire cdxi9006m = reg_1_4&cdxi5445m;
wire cdxi9007m = reg_1_3&cdxi6608m;
wire cdxi9008m = reg_1_2&cdxi5623m;
wire cdxi9009m = reg_1_1&cdxi5831m;
wire cdxi9010m = (cdxi8980m ^ cdxi8981m ^ cdxi8982m ^ cdxi8983m ^ cdxi8984m ^ cdxi8985m ^ cdxi8986m ^ cdxi8987m ^ cdxi8988m ^ cdxi8989m ^ cdxi8990m ^ cdxi8991m ^ cdxi8992m ^ cdxi8993m ^ cdxi8994m ^ cdxi8995m ^ cdxi8996m ^ cdxi8997m ^ cdxi8998m ^ cdxi8999m ^ cdxi9000m ^ cdxi9001m ^ cdxi9002m ^ cdxi9003m ^ cdxi9004m ^ cdxi9005m ^ cdxi9006m ^ cdxi9007m ^ cdxi9008m ^ cdxi9009m ^ cdxi7319m);
wire cdxi9011m = reg_1_0&cdxi9010m;
wire cdxi9012m = 0&0 ^ cdxi4711m ^ cdxi4722m ^ cdxi4762m ^ cdxi4732m;
wire cdxi9013m = a1&cdxi8562m;
wire cdxi9014m = reg_1_0&cdxi8566m;
wire cdxi9015m = a1&cdxi4810m;
wire cdxi9016m = reg_1_0&cdxi4815m;
wire cdxi9017m = cdxi4712m&cdxi4774m;
wire cdxi9018m = reg_1_1&cdxi4779m;
wire cdxi9019m = cdxi4743m&cdxi4955m;
wire cdxi9020m = cdxi5711m&r1m;
wire cdxi9021m = cdxi4875m&cdxi4763m;
wire cdxi9022m = cdxi4875m&cdxi4764m;
wire cdxi9023m = cdxi4953m&r7m;
wire cdxi9024m = cdxi4743m&cdxi4958m;
wire cdxi9025m = cdxi4743m&cdxi4959m;
wire cdxi9026m = cdxi4954m&r14m;
wire cdxi9027m = cdxi4916m&r15m;
wire cdxi9028m = cdxi4875m&r22m;
wire cdxi9029m = cdxi4762m&r29m;
wire cdxi9030m = cdxi4722m&r30m;
wire cdxi9031m = cdxi4743m&r37m;
wire cdxi9032m = cdxi4712m&r47m;
wire cdxi9033m = (cdxi67m ^ cdxi9019m ^ cdxi9020m ^ cdxi9021m ^ cdxi9022m ^ cdxi9023m ^ cdxi9024m ^ cdxi9025m ^ cdxi9026m ^ cdxi9027m ^ cdxi9028m ^ cdxi9029m ^ cdxi9030m ^ cdxi9031m ^ cdxi9032m);
wire cdxi9034m = a1&cdxi9033m;
wire cdxi9035m = reg_1_2&cdxi4965m;
wire cdxi9036m = reg_1_1&cdxi5039m;
wire cdxi9037m = reg_1_1&cdxi5040m;
wire cdxi9038m = reg_1_1&cdxi5041m;
wire cdxi9039m = reg_1_4&cdxi8875m;
wire cdxi9040m = reg_1_2&cdxi4968m;
wire cdxi9041m = reg_1_2&cdxi4969m;
wire cdxi9042m = reg_1_1&cdxi5042m;
wire cdxi9043m = reg_1_1&cdxi5043m;
wire cdxi9044m = reg_1_1&cdxi5044m;
wire cdxi9045m = reg_1_5&cdxi5331m;
wire cdxi9046m = reg_1_4&cdxi5368m;
wire cdxi9047m = reg_1_2&cdxi4964m;
wire cdxi9048m = reg_1_1&cdxi5038m;
wire cdxi9049m = (cdxi9035m ^ cdxi9036m ^ cdxi9037m ^ cdxi9038m ^ cdxi9039m ^ cdxi9040m ^ cdxi9041m ^ cdxi9042m ^ cdxi9043m ^ cdxi9044m ^ cdxi9045m ^ cdxi9046m ^ cdxi9047m ^ cdxi9048m ^ cdxi6261m);
wire cdxi9050m = reg_1_0&cdxi9049m;
wire cdxi9051m = cdxi4712m&cdxi5931m;
wire cdxi9052m = reg_1_1&cdxi5948m;
wire cdxi9053m = cdxi8487m;
wire cdxi9054m = 0&0 ^ a1 ^ cdxi4711m ^ cdxi4722m ^ cdxi4742m ^ cdxi4732m;
wire cdxi9055m = cdxi4742m&r0m;
wire cdxi9056m = cdxi4712m&r5m;
wire cdxi9057m = (cdxi11m ^ cdxi9055m ^ cdxi9056m);
wire cdxi9058m = a1&cdxi9057m;
wire cdxi9059m = reg_1_6&cdxi4664m;
wire cdxi9060m = reg_1_1&cdxi4689m;
wire cdxi9061m = (cdxi9059m ^ cdxi9060m ^ cdxi4905m);
wire cdxi9062m = reg_1_0&cdxi9061m;
wire cdxi9063m = 0&0 ^ a1 ^ cdxi4712m ^ cdxi4722m ^ cdxi4742m;
wire cdxi9064m = a1&cdxi5256m;
wire cdxi9065m = reg_1_0&cdxi5265m;
wire cdxi9066m = cdxi4743m&cdxi5143m;
wire cdxi9067m = reg_1_2&cdxi5152m;
wire cdxi9068m = cdxi4712m&cdxi5829m;
wire cdxi9069m = reg_1_1&cdxi5846m;







always @(posedge clk) begin
	reg_0_0 <= a0;
	reg_0_1 <= cdxi185m;
	reg_0_2 <= cdxi219m;
	reg_0_3 <= cdxi184m;
	reg_0_4 <= cdxi196m;
	reg_0_5 <= cdxi240m;
	reg_0_6 <= cdxi218m;
	reg_0_7 <= cdxi207m;
	reg_0_8 <= cdxi0m;
	reg_0_9 <= cdxi1m;
	reg_0_10 <= cdxi2m;
	reg_0_11 <= cdxi3m;
	reg_0_12 <= cdxi4m;
	reg_0_13 <= cdxi5m;
	reg_0_14 <= cdxi6m;
	reg_0_15 <= cdxi7m;
	reg_0_16 <= cdxi8m;
	reg_0_17 <= cdxi9m;
	reg_0_18 <= cdxi10m;
	reg_0_19 <= cdxi11m;
	reg_0_20 <= cdxi12m;
	reg_0_21 <= cdxi13m;
	reg_0_22 <= cdxi14m;
	reg_0_23 <= cdxi15m;
	reg_0_24 <= cdxi16m;
	reg_0_25 <= cdxi17m;
	reg_0_26 <= cdxi18m;
	reg_0_27 <= cdxi19m;
	reg_0_28 <= cdxi20m;
	reg_0_29 <= cdxi21m;
	reg_0_30 <= cdxi22m;
	reg_0_31 <= cdxi23m;
	reg_0_32 <= cdxi24m;
	reg_0_33 <= cdxi25m;
	reg_0_34 <= cdxi26m;
	reg_0_35 <= cdxi27m;
	reg_0_36 <= cdxi28m;
	reg_0_37 <= cdxi29m;
	reg_0_38 <= cdxi30m;
	reg_0_39 <= cdxi31m;
	reg_0_40 <= cdxi32m;
	reg_0_41 <= cdxi33m;
	reg_0_42 <= cdxi34m;
	reg_0_43 <= cdxi35m;
	reg_0_44 <= cdxi36m;
	reg_0_45 <= cdxi37m;
	reg_0_46 <= cdxi38m;
	reg_0_47 <= cdxi39m;
	reg_0_48 <= cdxi40m;
	reg_0_49 <= cdxi41m;
	reg_0_50 <= cdxi42m;
	reg_0_51 <= cdxi43m;
	reg_0_52 <= cdxi44m;
	reg_0_53 <= cdxi45m;
	reg_0_54 <= cdxi46m;
	reg_0_55 <= cdxi47m;
	reg_0_56 <= cdxi48m;
	reg_0_57 <= cdxi49m;
	reg_0_58 <= cdxi50m;
	reg_0_59 <= cdxi51m;
	reg_0_60 <= cdxi52m;
	reg_0_61 <= cdxi53m;
	reg_0_62 <= cdxi54m;
	reg_0_63 <= cdxi55m;
	reg_0_64 <= cdxi56m;
	reg_0_65 <= cdxi57m;
	reg_0_66 <= cdxi58m;
	reg_0_67 <= cdxi59m;
	reg_0_68 <= cdxi60m;
	reg_0_69 <= cdxi61m;
	reg_0_70 <= cdxi62m;
	reg_0_71 <= cdxi63m;
	reg_0_72 <= cdxi64m;
	reg_0_73 <= cdxi65m;
	reg_0_74 <= cdxi66m;
	reg_0_75 <= cdxi67m;
	reg_0_76 <= cdxi68m;
	reg_0_77 <= cdxi69m;
	reg_0_78 <= cdxi70m;
	reg_0_79 <= cdxi71m;
	reg_0_80 <= cdxi72m;
	reg_0_81 <= cdxi73m;
	reg_0_82 <= cdxi74m;
	reg_0_83 <= cdxi75m;
	reg_0_84 <= cdxi76m;
	reg_0_85 <= cdxi77m;
	reg_0_86 <= cdxi78m;
	reg_0_87 <= cdxi79m;
	reg_0_88 <= cdxi80m;
	reg_0_89 <= cdxi81m;
	reg_0_90 <= cdxi82m;
	reg_0_91 <= cdxi83m;
	reg_0_92 <= cdxi84m;
	reg_0_93 <= cdxi85m;
	reg_0_94 <= cdxi86m;
	reg_0_95 <= cdxi87m;
	reg_0_96 <= cdxi88m;
	reg_0_97 <= cdxi89m;
	reg_0_98 <= cdxi90m;
	reg_0_99 <= cdxi91m;
	reg_0_100 <= cdxi92m;
	reg_0_101 <= cdxi93m;
	reg_0_102 <= cdxi94m;
	reg_0_103 <= cdxi95m;
	reg_0_104 <= cdxi96m;
	reg_0_105 <= cdxi97m;
	reg_0_106 <= cdxi98m;
	reg_0_107 <= cdxi99m;
	reg_0_108 <= cdxi100m;
	reg_0_109 <= cdxi101m;
	reg_0_110 <= cdxi102m;
	reg_0_111 <= cdxi103m;
	reg_0_112 <= cdxi104m;
	reg_0_113 <= cdxi105m;
	reg_0_114 <= cdxi106m;
	reg_0_115 <= cdxi107m;
	reg_0_116 <= cdxi108m;
	reg_0_117 <= cdxi109m;
	reg_0_118 <= cdxi110m;
	reg_0_119 <= cdxi111m;
	reg_0_120 <= cdxi112m;
	reg_0_121 <= cdxi113m;
	reg_0_122 <= cdxi114m;
	reg_0_123 <= cdxi115m;
	reg_0_124 <= cdxi116m;
	reg_0_125 <= cdxi117m;
	reg_0_126 <= cdxi118m;
	reg_0_127 <= cdxi119m;
	reg_0_128 <= cdxi120m;
	reg_0_129 <= cdxi121m;
	reg_0_130 <= cdxi122m;
	reg_0_131 <= cdxi123m;
	reg_0_132 <= cdxi124m;
	reg_0_133 <= cdxi125m;
	reg_0_134 <= cdxi126m ^ cdxi129m ^ cdxi135m ^ cdxi141m ^ cdxi147m ^ cdxi153m ^ cdxi159m ^ cdxi163m ^ cdxi165m ^ cdxi169m ^ cdxi173m ^ cdxi175m ^ cdxi177m ^ cdxi179m ^ cdxi181m ^ cdxi189m ^ cdxi200m ^ cdxi211m ^ cdxi223m ^ cdxi233m ^ cdxi244m ^ cdxi254m ^ cdxi264m ^ cdxi274m ^ cdxi284m ^ cdxi294m ^ cdxi304m ^ cdxi314m ^ cdxi320m ^ cdxi322m ^ cdxi328m ^ cdxi334m ^ cdxi340m ^ cdxi346m ^ cdxi348m ^ cdxi350m ^ cdxi352m ^ cdxi354m ^ cdxi356m ^ cdxi358m ^ cdxi371m ^ cdxi393m ^ cdxi414m ^ cdxi434m ^ cdxi454m ^ cdxi474m ^ cdxi493m ^ cdxi512m ^ cdxi532m ^ cdxi551m ^ cdxi571m ^ cdxi590m ^ cdxi609m ^ cdxi627m ^ cdxi646m ^ cdxi665m ^ cdxi683m ^ cdxi701m ^ cdxi711m ^ cdxi713m ^ cdxi723m ^ cdxi741m ^ cdxi751m ^ cdxi753m ^ cdxi755m ^ cdxi765m ^ cdxi775m ^ cdxi785m ^ cdxi795m ^ cdxi797m ^ cdxi799m ^ cdxi809m ^ cdxi819m ^ cdxi841m ^ cdxi879m ^ cdxi918m ^ cdxi956m ^ cdxi994m ^ cdxi1030m ^ cdxi1067m ^ cdxi1104m ^ cdxi1140m ^ cdxi1177m ^ cdxi1212m ^ cdxi1249m ^ cdxi1284m ^ cdxi1320m ^ cdxi1355m ^ cdxi1390m ^ cdxi1426m ^ cdxi1460m ^ cdxi1495m ^ cdxi1529m ^ cdxi1564m ^ cdxi1598m ^ cdxi1616m ^ cdxi1634m ^ cdxi1668m ^ cdxi1702m ^ cdxi1720m ^ cdxi1722m ^ cdxi1724m ^ cdxi1742m ^ cdxi1797m ^ cdxi1869m ^ cdxi1938m ^ cdxi2009m ^ cdxi2078m ^ cdxi2149m ^ cdxi2219m ^ cdxi2288m ^ cdxi2357m ^ cdxi2424m ^ cdxi2492m ^ cdxi2560m ^ cdxi2626m ^ cdxi2693m ^ cdxi2727m ^ cdxi2729m ^ cdxi2763m ^ cdxi2797m ^ cdxi2870m ^ cdxi3008m ^ cdxi3143m ^ cdxi3277m ^ r126m;
	reg_0_135 <= cdxi3343m ^ cdxi141m ^ cdxi147m ^ cdxi153m ^ cdxi3344m ^ cdxi163m ^ cdxi169m ^ cdxi3346m ^ cdxi3348m ^ cdxi3350m ^ cdxi3352m ^ cdxi179m ^ cdxi3354m ^ cdxi3356m ^ cdxi3362m ^ cdxi200m ^ cdxi3371m ^ cdxi211m ^ cdxi3380m ^ cdxi3389m ^ cdxi223m ^ cdxi3394m ^ cdxi3396m ^ cdxi3398m ^ cdxi233m ^ cdxi244m ^ cdxi3400m ^ cdxi3402m ^ cdxi3404m ^ cdxi3406m ^ cdxi3408m ^ cdxi294m ^ cdxi3410m ^ cdxi3412m ^ cdxi314m ^ cdxi3414m ^ cdxi320m ^ cdxi3416m ^ cdxi3418m ^ cdxi346m ^ cdxi350m ^ cdxi352m ^ cdxi354m ^ cdxi356m ^ cdxi3420m ^ cdxi371m ^ cdxi3430m ^ cdxi393m ^ cdxi3447m ^ cdxi3464m ^ cdxi3481m ^ cdxi454m ^ cdxi474m ^ cdxi493m ^ cdxi512m ^ cdxi3490m ^ cdxi3500m ^ cdxi571m ^ cdxi3517m ^ cdxi609m ^ cdxi3526m ^ cdxi3536m ^ cdxi627m ^ cdxi3545m ^ cdxi3547m ^ cdxi683m ^ cdxi3549m ^ cdxi711m ^ cdxi741m ^ cdxi3551m ^ cdxi3553m ^ cdxi3555m ^ cdxi753m ^ cdxi765m ^ cdxi3557m ^ cdxi3559m ^ cdxi785m ^ cdxi3569m ^ cdxi3578m ^ cdxi797m ^ cdxi809m ^ cdxi3580m ^ cdxi3582m ^ cdxi841m ^ cdxi879m ^ cdxi994m ^ cdxi3600m ^ cdxi1030m ^ cdxi1140m ^ cdxi1177m ^ cdxi1249m ^ cdxi3633m ^ cdxi1390m ^ cdxi3666m ^ cdxi3699m ^ cdxi3716m ^ cdxi3718m ^ cdxi3720m ^ cdxi3722m ^ cdxi3724m ^ cdxi1616m ^ cdxi3726m ^ cdxi1634m ^ cdxi3728m ^ cdxi3730m ^ cdxi1702m ^ cdxi1720m ^ cdxi1724m ^ cdxi3732m ^ cdxi1797m ^ cdxi1869m ^ cdxi1938m ^ cdxi2009m ^ cdxi3766m ^ cdxi2078m ^ cdxi2219m ^ cdxi2357m ^ cdxi2424m ^ cdxi3831m ^ cdxi2492m ^ cdxi2763m ^ cdxi2797m ^ cdxi3931m ^ cdxi3277m ^ cdxi4639m ^ r127m;
	reg_0_136 <= cdxi4128m ^ cdxi129m ^ cdxi135m ^ cdxi141m ^ cdxi153m ^ cdxi163m ^ cdxi4129m ^ cdxi169m ^ cdxi4131m ^ cdxi4133m ^ cdxi177m ^ cdxi179m ^ cdxi181m ^ cdxi3362m ^ cdxi189m ^ cdxi211m ^ cdxi3389m ^ cdxi3394m ^ cdxi3396m ^ cdxi233m ^ cdxi3400m ^ cdxi3402m ^ cdxi264m ^ cdxi4139m ^ cdxi4144m ^ cdxi4146m ^ cdxi294m ^ cdxi3410m ^ cdxi4148m ^ cdxi4150m ^ cdxi3412m ^ cdxi314m ^ cdxi3416m ^ cdxi334m ^ cdxi3418m ^ cdxi340m ^ cdxi346m ^ cdxi348m ^ cdxi352m ^ cdxi4152m ^ cdxi3420m ^ cdxi371m ^ cdxi3464m ^ cdxi474m ^ cdxi4162m ^ cdxi493m ^ cdxi4179m ^ cdxi4188m ^ cdxi3490m ^ cdxi3500m ^ cdxi4190m ^ cdxi590m ^ cdxi609m ^ cdxi3536m ^ cdxi627m ^ cdxi646m ^ cdxi3545m ^ cdxi3547m ^ cdxi3549m ^ cdxi711m ^ cdxi723m ^ cdxi741m ^ cdxi3553m ^ cdxi753m ^ cdxi4192m ^ cdxi755m ^ cdxi4194m ^ cdxi3557m ^ cdxi3569m ^ cdxi799m ^ cdxi3580m ^ cdxi3582m ^ cdxi841m ^ cdxi918m ^ cdxi3600m ^ cdxi1067m ^ cdxi1104m ^ cdxi1140m ^ cdxi4212m ^ cdxi1249m ^ cdxi1284m ^ cdxi3633m ^ cdxi1320m ^ cdxi1426m ^ cdxi1529m ^ cdxi3699m ^ cdxi4229m ^ cdxi1564m ^ cdxi3720m ^ cdxi1598m ^ cdxi4231m ^ cdxi4233m ^ cdxi3726m ^ cdxi4235m ^ cdxi1668m ^ cdxi3730m ^ cdxi1720m ^ cdxi1722m ^ cdxi1724m ^ cdxi2009m ^ cdxi2149m ^ cdxi2219m ^ cdxi2288m ^ cdxi4269m ^ cdxi4302m ^ cdxi4304m ^ cdxi4370m ^ cdxi3143m ^ cdxi4639m ^ cdxi4436m ^ r128m;
	reg_0_137 <= cdxi4438m ^ cdxi129m ^ cdxi135m ^ cdxi141m ^ cdxi153m ^ cdxi4129m ^ cdxi165m ^ cdxi169m ^ cdxi3346m ^ cdxi3348m ^ cdxi173m ^ cdxi175m ^ cdxi177m ^ cdxi181m ^ cdxi3354m ^ cdxi3356m ^ cdxi3362m ^ cdxi189m ^ cdxi200m ^ cdxi3371m ^ cdxi211m ^ cdxi3394m ^ cdxi233m ^ cdxi3400m ^ cdxi3402m ^ cdxi254m ^ cdxi4139m ^ cdxi3406m ^ cdxi4144m ^ cdxi274m ^ cdxi284m ^ cdxi4146m ^ cdxi294m ^ cdxi4439m ^ cdxi4441m ^ cdxi3412m ^ cdxi3414m ^ cdxi334m ^ cdxi348m ^ cdxi354m ^ cdxi4443m ^ cdxi358m ^ cdxi4453m ^ cdxi393m ^ cdxi3481m ^ cdxi4162m ^ cdxi512m ^ cdxi3490m ^ cdxi532m ^ cdxi551m ^ cdxi571m ^ cdxi4190m ^ cdxi3517m ^ cdxi627m ^ cdxi646m ^ cdxi665m ^ cdxi3547m ^ cdxi683m ^ cdxi3549m ^ cdxi713m ^ cdxi741m ^ cdxi4192m ^ cdxi755m ^ cdxi4194m ^ cdxi765m ^ cdxi3557m ^ cdxi3559m ^ cdxi797m ^ cdxi799m ^ cdxi819m ^ cdxi841m ^ cdxi879m ^ cdxi918m ^ cdxi956m ^ cdxi994m ^ cdxi4478m ^ cdxi4511m ^ cdxi1104m ^ cdxi4528m ^ cdxi1355m ^ cdxi1390m ^ cdxi1426m ^ cdxi4530m ^ cdxi3718m ^ cdxi3720m ^ cdxi3722m ^ cdxi3724m ^ cdxi1616m ^ cdxi4235m ^ cdxi1634m ^ cdxi3730m ^ cdxi1702m ^ cdxi1720m ^ cdxi1724m ^ cdxi3732m ^ cdxi1742m ^ cdxi1797m ^ cdxi4564m ^ cdxi2009m ^ cdxi2078m ^ cdxi2149m ^ cdxi2219m ^ cdxi2288m ^ cdxi4269m ^ cdxi3831m ^ cdxi2492m ^ cdxi2626m ^ cdxi2693m ^ cdxi2727m ^ cdxi2763m ^ cdxi4302m ^ cdxi2797m ^ cdxi4304m ^ cdxi4370m ^ cdxi3143m ^ cdxi3277m ^ r129m;
	reg_0_138 <= cdxi4597m ^ cdxi129m ^ cdxi135m ^ cdxi3344m ^ cdxi4129m ^ cdxi165m ^ cdxi169m ^ cdxi3348m ^ cdxi4131m ^ cdxi3350m ^ cdxi179m ^ cdxi181m ^ cdxi3362m ^ cdxi189m ^ cdxi200m ^ cdxi211m ^ cdxi4598m ^ cdxi3380m ^ cdxi223m ^ cdxi4600m ^ cdxi233m ^ cdxi244m ^ cdxi3400m ^ cdxi3404m ^ cdxi4139m ^ cdxi3406m ^ cdxi3408m ^ cdxi4144m ^ cdxi274m ^ cdxi284m ^ cdxi294m ^ cdxi4439m ^ cdxi4441m ^ cdxi3410m ^ cdxi4602m ^ cdxi4148m ^ cdxi4150m ^ cdxi3412m ^ cdxi314m ^ cdxi320m ^ cdxi3416m ^ cdxi334m ^ cdxi3418m ^ cdxi352m ^ cdxi354m ^ cdxi4443m ^ cdxi356m ^ cdxi4152m ^ cdxi3430m ^ cdxi4453m ^ cdxi3447m ^ cdxi414m ^ cdxi3464m ^ cdxi3500m ^ cdxi532m ^ cdxi551m ^ cdxi571m ^ cdxi3517m ^ cdxi590m ^ cdxi609m ^ cdxi3526m ^ cdxi646m ^ cdxi3545m ^ cdxi3547m ^ cdxi713m ^ cdxi741m ^ cdxi3551m ^ cdxi751m ^ cdxi3555m ^ cdxi753m ^ cdxi4194m ^ cdxi797m ^ cdxi809m ^ cdxi3582m ^ cdxi841m ^ cdxi918m ^ cdxi4620m ^ cdxi994m ^ cdxi3600m ^ cdxi1030m ^ cdxi4478m ^ cdxi1067m ^ cdxi1212m ^ cdxi1284m ^ cdxi1355m ^ cdxi1390m ^ cdxi1460m ^ cdxi1495m ^ cdxi1529m ^ cdxi3699m ^ cdxi1564m ^ cdxi3720m ^ cdxi3722m ^ cdxi4637m ^ cdxi4231m ^ cdxi1616m ^ cdxi4233m ^ cdxi4235m ^ cdxi3730m ^ cdxi1702m ^ cdxi1724m ^ cdxi3732m ^ cdxi1797m ^ cdxi1869m ^ cdxi4564m ^ cdxi1938m ^ cdxi2009m ^ cdxi2149m ^ cdxi2288m ^ cdxi4269m ^ cdxi2626m ^ cdxi2693m ^ cdxi2727m ^ cdxi4302m ^ cdxi2797m ^ cdxi2870m ^ cdxi3008m ^ cdxi4639m ^ r130m;
	reg_0_139 <= cdxi129m ^ cdxi147m ^ cdxi153m ^ cdxi159m ^ cdxi3344m ^ cdxi4129m ^ cdxi165m ^ cdxi169m ^ cdxi3346m ^ cdxi3348m ^ cdxi175m ^ cdxi3352m ^ cdxi179m ^ cdxi181m ^ cdxi3354m ^ cdxi3356m ^ cdxi211m ^ cdxi4598m ^ cdxi3380m ^ cdxi3389m ^ cdxi223m ^ cdxi3394m ^ cdxi3396m ^ cdxi4600m ^ cdxi233m ^ cdxi3402m ^ cdxi4139m ^ cdxi3408m ^ cdxi294m ^ cdxi4602m ^ cdxi4148m ^ cdxi3412m ^ cdxi314m ^ cdxi3414m ^ cdxi3416m ^ cdxi334m ^ cdxi3418m ^ cdxi340m ^ cdxi346m ^ cdxi348m ^ cdxi352m ^ cdxi354m ^ cdxi4443m ^ cdxi358m ^ cdxi371m ^ cdxi3447m ^ cdxi3464m ^ cdxi434m ^ cdxi454m ^ cdxi4162m ^ cdxi493m ^ cdxi512m ^ cdxi3490m ^ cdxi3500m ^ cdxi532m ^ cdxi3526m ^ cdxi3545m ^ cdxi665m ^ cdxi3547m ^ cdxi683m ^ cdxi723m ^ cdxi741m ^ cdxi3551m ^ cdxi751m ^ cdxi3553m ^ cdxi753m ^ cdxi4192m ^ cdxi755m ^ cdxi4194m ^ cdxi3557m ^ cdxi775m ^ cdxi3559m ^ cdxi3569m ^ cdxi797m ^ cdxi809m ^ cdxi819m ^ cdxi3582m ^ cdxi841m ^ cdxi879m ^ cdxi956m ^ cdxi4620m ^ cdxi994m ^ cdxi3600m ^ cdxi1030m ^ cdxi1067m ^ cdxi4511m ^ cdxi1104m ^ cdxi1177m ^ cdxi1212m ^ cdxi1284m ^ cdxi3633m ^ cdxi1355m ^ cdxi1390m ^ cdxi1460m ^ cdxi3666m ^ cdxi3716m ^ cdxi1564m ^ cdxi3718m ^ cdxi3724m ^ cdxi4637m ^ cdxi4231m ^ cdxi1616m ^ cdxi3726m ^ cdxi4235m ^ cdxi3728m ^ cdxi1720m ^ cdxi3732m ^ cdxi1742m ^ cdxi1869m ^ cdxi4564m ^ cdxi1938m ^ cdxi2078m ^ cdxi2149m ^ cdxi2219m ^ cdxi2357m ^ cdxi4269m ^ cdxi3831m ^ cdxi2727m ^ cdxi4302m ^ cdxi2797m ^ cdxi4304m ^ cdxi3931m ^ cdxi3008m ^ cdxi3277m ^ cdxi4639m ^ r131m;
	reg_0_140 <= cdxi4640m ^ cdxi153m ^ cdxi3344m ^ cdxi169m ^ cdxi3348m ^ cdxi4131m ^ cdxi3350m ^ cdxi3352m ^ cdxi179m ^ cdxi181m ^ cdxi3356m ^ cdxi200m ^ cdxi4645m ^ cdxi211m ^ cdxi223m ^ cdxi3394m ^ cdxi4600m ^ cdxi244m ^ cdxi3402m ^ cdxi264m ^ cdxi3404m ^ cdxi4139m ^ cdxi3408m ^ cdxi274m ^ cdxi284m ^ cdxi4146m ^ cdxi4439m ^ cdxi4602m ^ cdxi3412m ^ cdxi314m ^ cdxi322m ^ cdxi340m ^ cdxi348m ^ cdxi4443m ^ cdxi356m ^ cdxi358m ^ cdxi371m ^ cdxi3447m ^ cdxi414m ^ cdxi3464m ^ cdxi3481m ^ cdxi4162m ^ cdxi493m ^ cdxi4179m ^ cdxi512m ^ cdxi3500m ^ cdxi571m ^ cdxi3517m ^ cdxi590m ^ cdxi3526m ^ cdxi627m ^ cdxi711m ^ cdxi713m ^ cdxi741m ^ cdxi3551m ^ cdxi3553m ^ cdxi753m ^ cdxi765m ^ cdxi3569m ^ cdxi819m ^ cdxi3580m ^ cdxi3582m ^ cdxi841m ^ cdxi879m ^ cdxi918m ^ cdxi956m ^ cdxi994m ^ cdxi3600m ^ cdxi1030m ^ cdxi4478m ^ cdxi1067m ^ cdxi4511m ^ cdxi1177m ^ cdxi4212m ^ cdxi1249m ^ cdxi1320m ^ cdxi1355m ^ cdxi1390m ^ cdxi1426m ^ cdxi1460m ^ cdxi1495m ^ cdxi1529m ^ cdxi3666m ^ cdxi4530m ^ cdxi1564m ^ cdxi3718m ^ cdxi3720m ^ cdxi3722m ^ cdxi4637m ^ cdxi1616m ^ cdxi4233m ^ cdxi3726m ^ cdxi4235m ^ cdxi1634m ^ cdxi3728m ^ cdxi1720m ^ cdxi1722m ^ cdxi1869m ^ cdxi3766m ^ cdxi2078m ^ cdxi2492m ^ cdxi2560m ^ cdxi2626m ^ cdxi2763m ^ cdxi4304m ^ cdxi3931m ^ cdxi4639m ^ cdxi4436m ^ r132m;
	reg_0_141 <= cdxi4650m ^ cdxi129m ^ cdxi153m ^ cdxi3344m ^ cdxi165m ^ cdxi3346m ^ cdxi3348m ^ cdxi3350m ^ cdxi179m ^ cdxi181m ^ cdxi3362m ^ cdxi189m ^ cdxi3371m ^ cdxi211m ^ cdxi4598m ^ cdxi3380m ^ cdxi3394m ^ cdxi3398m ^ cdxi4600m ^ cdxi233m ^ cdxi244m ^ cdxi4139m ^ cdxi284m ^ cdxi4146m ^ cdxi294m ^ cdxi304m ^ cdxi3410m ^ cdxi4602m ^ cdxi4150m ^ cdxi314m ^ cdxi320m ^ cdxi3416m ^ cdxi322m ^ cdxi334m ^ cdxi340m ^ cdxi348m ^ cdxi350m ^ cdxi354m ^ cdxi358m ^ cdxi3420m ^ cdxi371m ^ cdxi3481m ^ cdxi434m ^ cdxi474m ^ cdxi4162m ^ cdxi4179m ^ cdxi3490m ^ cdxi3517m ^ cdxi590m ^ cdxi609m ^ cdxi646m ^ cdxi3545m ^ cdxi4651m ^ cdxi665m ^ cdxi3547m ^ cdxi713m ^ cdxi741m ^ cdxi3551m ^ cdxi751m ^ cdxi3553m ^ cdxi4192m ^ cdxi755m ^ cdxi3559m ^ cdxi4653m ^ cdxi797m ^ cdxi3580m ^ cdxi3582m ^ cdxi841m ^ cdxi956m ^ cdxi4620m ^ cdxi994m ^ cdxi3600m ^ cdxi1030m ^ cdxi4478m ^ cdxi4511m ^ cdxi1177m ^ cdxi4212m ^ cdxi1320m ^ cdxi4528m ^ cdxi1426m ^ cdxi1460m ^ cdxi1495m ^ cdxi3666m ^ cdxi3699m ^ cdxi4229m ^ cdxi3720m ^ cdxi1598m ^ cdxi4655m ^ cdxi3724m ^ cdxi4637m ^ cdxi4231m ^ cdxi1616m ^ cdxi3726m ^ cdxi4235m ^ cdxi3728m ^ cdxi3730m ^ cdxi1702m ^ cdxi1724m ^ cdxi1742m ^ cdxi1797m ^ cdxi1938m ^ cdxi2009m ^ cdxi2219m ^ cdxi2288m ^ cdxi3831m ^ cdxi2492m ^ cdxi2626m ^ cdxi2693m ^ cdxi2727m ^ cdxi2797m ^ cdxi4304m ^ cdxi3931m ^ cdxi3008m ^ cdxi4639m ^ r133m;





	reg_1_0 <= a1;
	reg_1_1 <= cdxi4712m;
	reg_1_2 <= cdxi4743m;
	reg_1_3 <= cdxi4711m;
	reg_1_4 <= cdxi4722m;
	reg_1_5 <= cdxi4762m;
	reg_1_6 <= cdxi4742m;
	reg_1_7 <= cdxi4732m;
	reg_1_8 <= cdxi128m;
	reg_1_9 <= cdxi134m;
	reg_1_10 <= cdxi140m;
	reg_1_11 <= cdxi146m;
	reg_1_12 <= cdxi152m;
	reg_1_13 <= cdxi158m;
	reg_1_14 <= cdxi168m;
	reg_1_15 <= cdxi3358m;
	reg_1_16 <= cdxi183m;
	reg_1_17 <= cdxi195m;
	reg_1_18 <= cdxi3367m;
	reg_1_19 <= cdxi4641m;
	reg_1_20 <= cdxi206m;
	reg_1_21 <= cdxi4135m;
	reg_1_22 <= cdxi3376m;
	reg_1_23 <= cdxi3385m;
	reg_1_24 <= cdxi217m;
	reg_1_25 <= cdxi270m;
	reg_1_26 <= cdxi280m;
	reg_1_27 <= cdxi310m;
	reg_1_28 <= cdxi290m;
	reg_1_29 <= cdxi229m;
	reg_1_30 <= cdxi239m;
	reg_1_31 <= cdxi300m;
	reg_1_32 <= cdxi324m;
	reg_1_33 <= cdxi250m;
	reg_1_34 <= cdxi260m;
	reg_1_35 <= cdxi336m;
	reg_1_36 <= cdxi360m;
	reg_1_37 <= cdxi3422m;
	reg_1_38 <= cdxi4445m;
	reg_1_39 <= cdxi383m;
	reg_1_40 <= cdxi3439m;
	reg_1_41 <= cdxi404m;
	reg_1_42 <= cdxi3456m;
	reg_1_43 <= cdxi3473m;
	reg_1_44 <= cdxi424m;
	reg_1_45 <= cdxi444m;
	reg_1_46 <= cdxi465m;
	reg_1_47 <= cdxi4657m;
	reg_1_48 <= cdxi4154m;
	reg_1_49 <= cdxi484m;
	reg_1_50 <= cdxi4171m;
	reg_1_51 <= cdxi503m;
	reg_1_52 <= cdxi675m;
	reg_1_53 <= cdxi693m;
	reg_1_54 <= cdxi3492m;
	reg_1_55 <= cdxi523m;
	reg_1_56 <= cdxi543m;
	reg_1_57 <= cdxi561m;
	reg_1_58 <= cdxi715m;
	reg_1_59 <= cdxi733m;
	reg_1_60 <= cdxi3509m;
	reg_1_61 <= cdxi581m;
	reg_1_62 <= cdxi600m;
	reg_1_63 <= cdxi777m;
	reg_1_64 <= cdxi3528m;
	reg_1_65 <= cdxi619m;
	reg_1_66 <= cdxi3561m;
	reg_1_67 <= cdxi637m;
	reg_1_68 <= cdxi801m;
	reg_1_69 <= cdxi757m;
	reg_1_70 <= cdxi656m;
	reg_1_71 <= cdxi821m;
	reg_1_72 <= cdxi860m;
	reg_1_73 <= cdxi899m;
	reg_1_74 <= cdxi937m;
	reg_1_75 <= cdxi4604m;
	reg_1_76 <= cdxi976m;
	reg_1_77 <= cdxi3584m;
	reg_1_78 <= cdxi1012m;
	reg_1_79 <= cdxi4462m;
	reg_1_80 <= cdxi1049m;
	reg_1_81 <= cdxi4495m;
	reg_1_82 <= cdxi1087m;
	reg_1_83 <= cdxi1122m;
	reg_1_84 <= cdxi4658m;
	reg_1_85 <= cdxi1159m;
	reg_1_86 <= cdxi1195m;
	reg_1_87 <= cdxi4196m;
	reg_1_88 <= cdxi1231m;
	reg_1_89 <= cdxi1267m;
	reg_1_90 <= cdxi3617m;
	reg_1_91 <= cdxi1302m;
	reg_1_92 <= cdxi1582m;
	reg_1_93 <= cdxi1338m;
	reg_1_94 <= cdxi1373m;
	reg_1_95 <= cdxi1409m;
	reg_1_96 <= cdxi1444m;
	reg_1_97 <= cdxi1478m;
	reg_1_98 <= cdxi1513m;
	reg_1_99 <= cdxi3650m;
	reg_1_100 <= cdxi3683m;
	reg_1_101 <= cdxi1686m;
	reg_1_102 <= cdxi1618m;
	reg_1_103 <= cdxi1652m;
	reg_1_104 <= cdxi1547m;
	reg_1_105 <= cdxi1726m;
	reg_1_106 <= cdxi1760m;
	reg_1_107 <= cdxi1833m;
	reg_1_108 <= cdxi4532m;
	reg_1_109 <= cdxi1903m;
	reg_1_110 <= cdxi1973m;
	reg_1_111 <= cdxi3734m;
	reg_1_112 <= cdxi2044m;
	reg_1_113 <= cdxi4659m;
	reg_1_114 <= cdxi2113m;
	reg_1_115 <= cdxi2185m;
	reg_1_116 <= cdxi2255m;
	reg_1_117 <= cdxi2322m;
	reg_1_118 <= cdxi4660m;
	reg_1_119 <= cdxi4237m;
	reg_1_120 <= cdxi2391m;
	reg_1_121 <= cdxi3799m;
	reg_1_122 <= cdxi2458m;
	reg_1_123 <= cdxi2526m;
	reg_1_124 <= cdxi2731m;
	reg_1_125 <= cdxi2594m;
	reg_1_126 <= cdxi2660m;
	reg_1_127 <= cdxi3865m;
	reg_1_128 <= cdxi4306m;
	reg_1_129 <= cdxi2799m;
	reg_1_130 <= cdxi2939m;
	reg_1_131 <= cdxi3075m;
	reg_1_132 <= cdxi3210m;
	reg_1_133 <= cdxi3997m;
	reg_1_134 <= cdxi4661m ^ cdxi4663m ^ cdxi4668m ^ cdxi4673m ^ cdxi4678m ^ cdxi4683m ^ cdxi4688m ^ cdxi4692m ^ cdxi4694m ^ cdxi4697m ^ cdxi4701m ^ cdxi4703m ^ cdxi4705m ^ cdxi4707m ^ cdxi4709m ^ cdxi4716m ^ cdxi4726m ^ cdxi4736m ^ cdxi4747m ^ cdxi4756m ^ cdxi4766m ^ cdxi4775m ^ cdxi4784m ^ cdxi4793m ^ cdxi4802m ^ cdxi4811m ^ cdxi4820m ^ cdxi4829m ^ cdxi4835m ^ cdxi4837m ^ cdxi4842m ^ cdxi4848m ^ cdxi4853m ^ cdxi4859m ^ cdxi4861m ^ cdxi4863m ^ cdxi4865m ^ cdxi4867m ^ cdxi4869m ^ cdxi4871m ^ cdxi4883m ^ cdxi4904m ^ cdxi4924m ^ cdxi4943m ^ cdxi4962m ^ cdxi4981m ^ cdxi4999m ^ cdxi5017m ^ cdxi5036m ^ cdxi5054m ^ cdxi5073m ^ cdxi5091m ^ cdxi5109m ^ cdxi5126m ^ cdxi5144m ^ cdxi5162m ^ cdxi5179m ^ cdxi5196m ^ cdxi5206m ^ cdxi5208m ^ cdxi5217m ^ cdxi5234m ^ cdxi5244m ^ cdxi5246m ^ cdxi5248m ^ cdxi5257m ^ cdxi5267m ^ cdxi5276m ^ cdxi5286m ^ cdxi5288m ^ cdxi5290m ^ cdxi5299m ^ cdxi5309m ^ cdxi5330m ^ cdxi5367m ^ cdxi5405m ^ cdxi5442m ^ cdxi5479m ^ cdxi5514m ^ cdxi5550m ^ cdxi5586m ^ cdxi5621m ^ cdxi5657m ^ cdxi5691m ^ cdxi5727m ^ cdxi5761m ^ cdxi5796m ^ cdxi5830m ^ cdxi5864m ^ cdxi5899m ^ cdxi5932m ^ cdxi5966m ^ cdxi5999m ^ cdxi6033m ^ cdxi6066m ^ cdxi6084m ^ cdxi6101m ^ cdxi6134m ^ cdxi6167m ^ cdxi6185m ^ cdxi6187m ^ cdxi6189m ^ cdxi6206m ^ cdxi6260m ^ cdxi6331m ^ cdxi6399m ^ cdxi6469m ^ cdxi6537m ^ cdxi6607m ^ cdxi6676m ^ cdxi6744m ^ cdxi6812m ^ cdxi6878m ^ cdxi6945m ^ cdxi7012m ^ cdxi7077m ^ cdxi7143m ^ cdxi7177m ^ cdxi7179m ^ cdxi7212m ^ cdxi7246m ^ cdxi7318m ^ cdxi7455m ^ cdxi7589m ^ cdxi7722m ^ r126m;
	reg_1_135 <= cdxi7788m ^ cdxi4673m ^ cdxi4678m ^ cdxi4683m ^ cdxi7789m ^ cdxi4692m ^ cdxi4697m ^ cdxi7791m ^ cdxi7793m ^ cdxi7795m ^ cdxi7797m ^ cdxi4707m ^ cdxi7799m ^ cdxi7801m ^ cdxi7806m ^ cdxi4726m ^ cdxi7814m ^ cdxi4736m ^ cdxi7822m ^ cdxi7830m ^ cdxi4747m ^ cdxi7835m ^ cdxi7837m ^ cdxi7839m ^ cdxi4756m ^ cdxi4766m ^ cdxi7841m ^ cdxi7843m ^ cdxi7845m ^ cdxi7847m ^ cdxi7849m ^ cdxi4811m ^ cdxi7851m ^ cdxi7853m ^ cdxi4829m ^ cdxi7855m ^ cdxi4835m ^ cdxi7857m ^ cdxi7859m ^ cdxi4859m ^ cdxi4863m ^ cdxi4865m ^ cdxi4867m ^ cdxi4869m ^ cdxi7861m ^ cdxi4883m ^ cdxi7870m ^ cdxi4904m ^ cdxi7886m ^ cdxi7902m ^ cdxi7918m ^ cdxi4962m ^ cdxi4981m ^ cdxi4999m ^ cdxi5017m ^ cdxi7927m ^ cdxi7936m ^ cdxi5073m ^ cdxi7952m ^ cdxi5109m ^ cdxi7961m ^ cdxi7970m ^ cdxi5126m ^ cdxi7979m ^ cdxi7981m ^ cdxi5179m ^ cdxi7983m ^ cdxi5206m ^ cdxi5234m ^ cdxi7985m ^ cdxi7987m ^ cdxi7989m ^ cdxi5246m ^ cdxi5257m ^ cdxi7991m ^ cdxi7993m ^ cdxi5276m ^ cdxi8002m ^ cdxi8011m ^ cdxi5288m ^ cdxi5299m ^ cdxi8013m ^ cdxi8015m ^ cdxi5330m ^ cdxi5367m ^ cdxi5479m ^ cdxi8032m ^ cdxi5514m ^ cdxi5621m ^ cdxi5657m ^ cdxi5727m ^ cdxi8064m ^ cdxi5864m ^ cdxi8096m ^ cdxi8128m ^ cdxi8145m ^ cdxi8147m ^ cdxi8149m ^ cdxi8151m ^ cdxi8153m ^ cdxi6084m ^ cdxi8155m ^ cdxi6101m ^ cdxi8157m ^ cdxi8159m ^ cdxi6167m ^ cdxi6185m ^ cdxi6189m ^ cdxi8161m ^ cdxi6260m ^ cdxi6331m ^ cdxi6399m ^ cdxi6469m ^ cdxi8194m ^ cdxi6537m ^ cdxi6676m ^ cdxi6812m ^ cdxi6878m ^ cdxi8258m ^ cdxi6945m ^ cdxi7212m ^ cdxi7246m ^ cdxi8357m ^ cdxi7722m ^ cdxi9053m ^ r127m;
	reg_1_136 <= cdxi8553m ^ cdxi4663m ^ cdxi4668m ^ cdxi4673m ^ cdxi4683m ^ cdxi4692m ^ cdxi8554m ^ cdxi4697m ^ cdxi8556m ^ cdxi8558m ^ cdxi4705m ^ cdxi4707m ^ cdxi4709m ^ cdxi7806m ^ cdxi4716m ^ cdxi4736m ^ cdxi7830m ^ cdxi7835m ^ cdxi7837m ^ cdxi4756m ^ cdxi7841m ^ cdxi7843m ^ cdxi4784m ^ cdxi8563m ^ cdxi8568m ^ cdxi8570m ^ cdxi4811m ^ cdxi7851m ^ cdxi8572m ^ cdxi8574m ^ cdxi7853m ^ cdxi4829m ^ cdxi7857m ^ cdxi4848m ^ cdxi7859m ^ cdxi4853m ^ cdxi4859m ^ cdxi4861m ^ cdxi4865m ^ cdxi8576m ^ cdxi7861m ^ cdxi4883m ^ cdxi7902m ^ cdxi4981m ^ cdxi8585m ^ cdxi4999m ^ cdxi8601m ^ cdxi8610m ^ cdxi7927m ^ cdxi7936m ^ cdxi8612m ^ cdxi5091m ^ cdxi5109m ^ cdxi7970m ^ cdxi5126m ^ cdxi5144m ^ cdxi7979m ^ cdxi7981m ^ cdxi7983m ^ cdxi5206m ^ cdxi5217m ^ cdxi5234m ^ cdxi7987m ^ cdxi5246m ^ cdxi8614m ^ cdxi5248m ^ cdxi8616m ^ cdxi7991m ^ cdxi8002m ^ cdxi5290m ^ cdxi8013m ^ cdxi8015m ^ cdxi5330m ^ cdxi5405m ^ cdxi8032m ^ cdxi5550m ^ cdxi5586m ^ cdxi5621m ^ cdxi8633m ^ cdxi5727m ^ cdxi5761m ^ cdxi8064m ^ cdxi5796m ^ cdxi5899m ^ cdxi5999m ^ cdxi8128m ^ cdxi8650m ^ cdxi6033m ^ cdxi8149m ^ cdxi6066m ^ cdxi8652m ^ cdxi8654m ^ cdxi8155m ^ cdxi8656m ^ cdxi6134m ^ cdxi8159m ^ cdxi6185m ^ cdxi6187m ^ cdxi6189m ^ cdxi6469m ^ cdxi6607m ^ cdxi6676m ^ cdxi6744m ^ cdxi8689m ^ cdxi8722m ^ cdxi8724m ^ cdxi8789m ^ cdxi7589m ^ cdxi9053m ^ cdxi8855m ^ r128m;
	reg_1_137 <= cdxi8857m ^ cdxi4663m ^ cdxi4668m ^ cdxi4673m ^ cdxi4683m ^ cdxi8554m ^ cdxi4694m ^ cdxi4697m ^ cdxi7791m ^ cdxi7793m ^ cdxi4701m ^ cdxi4703m ^ cdxi4705m ^ cdxi4709m ^ cdxi7799m ^ cdxi7801m ^ cdxi7806m ^ cdxi4716m ^ cdxi4726m ^ cdxi7814m ^ cdxi4736m ^ cdxi7835m ^ cdxi4756m ^ cdxi7841m ^ cdxi7843m ^ cdxi4775m ^ cdxi8563m ^ cdxi7847m ^ cdxi8568m ^ cdxi4793m ^ cdxi4802m ^ cdxi8570m ^ cdxi4811m ^ cdxi8858m ^ cdxi8860m ^ cdxi7853m ^ cdxi7855m ^ cdxi4848m ^ cdxi4861m ^ cdxi4867m ^ cdxi8862m ^ cdxi4871m ^ cdxi8871m ^ cdxi4904m ^ cdxi7918m ^ cdxi8585m ^ cdxi5017m ^ cdxi7927m ^ cdxi5036m ^ cdxi5054m ^ cdxi5073m ^ cdxi8612m ^ cdxi7952m ^ cdxi5126m ^ cdxi5144m ^ cdxi5162m ^ cdxi7981m ^ cdxi5179m ^ cdxi7983m ^ cdxi5208m ^ cdxi5234m ^ cdxi8614m ^ cdxi5248m ^ cdxi8616m ^ cdxi5257m ^ cdxi7991m ^ cdxi7993m ^ cdxi5288m ^ cdxi5290m ^ cdxi5309m ^ cdxi5330m ^ cdxi5367m ^ cdxi5405m ^ cdxi5442m ^ cdxi5479m ^ cdxi8895m ^ cdxi8927m ^ cdxi5586m ^ cdxi8944m ^ cdxi5830m ^ cdxi5864m ^ cdxi5899m ^ cdxi8946m ^ cdxi8147m ^ cdxi8149m ^ cdxi8151m ^ cdxi8153m ^ cdxi6084m ^ cdxi8656m ^ cdxi6101m ^ cdxi8159m ^ cdxi6167m ^ cdxi6185m ^ cdxi6189m ^ cdxi8161m ^ cdxi6206m ^ cdxi6260m ^ cdxi8979m ^ cdxi6469m ^ cdxi6537m ^ cdxi6607m ^ cdxi6676m ^ cdxi6744m ^ cdxi8689m ^ cdxi8258m ^ cdxi6945m ^ cdxi7077m ^ cdxi7143m ^ cdxi7177m ^ cdxi7212m ^ cdxi8722m ^ cdxi7246m ^ cdxi8724m ^ cdxi8789m ^ cdxi7589m ^ cdxi7722m ^ r129m;
	reg_1_138 <= cdxi9012m ^ cdxi4663m ^ cdxi4668m ^ cdxi7789m ^ cdxi8554m ^ cdxi4694m ^ cdxi4697m ^ cdxi7793m ^ cdxi8556m ^ cdxi7795m ^ cdxi4707m ^ cdxi4709m ^ cdxi7806m ^ cdxi4716m ^ cdxi4726m ^ cdxi4736m ^ cdxi9013m ^ cdxi7822m ^ cdxi4747m ^ cdxi9015m ^ cdxi4756m ^ cdxi4766m ^ cdxi7841m ^ cdxi7845m ^ cdxi8563m ^ cdxi7847m ^ cdxi7849m ^ cdxi8568m ^ cdxi4793m ^ cdxi4802m ^ cdxi4811m ^ cdxi8858m ^ cdxi8860m ^ cdxi7851m ^ cdxi9017m ^ cdxi8572m ^ cdxi8574m ^ cdxi7853m ^ cdxi4829m ^ cdxi4835m ^ cdxi7857m ^ cdxi4848m ^ cdxi7859m ^ cdxi4865m ^ cdxi4867m ^ cdxi8862m ^ cdxi4869m ^ cdxi8576m ^ cdxi7870m ^ cdxi8871m ^ cdxi7886m ^ cdxi4924m ^ cdxi7902m ^ cdxi7936m ^ cdxi5036m ^ cdxi5054m ^ cdxi5073m ^ cdxi7952m ^ cdxi5091m ^ cdxi5109m ^ cdxi7961m ^ cdxi5144m ^ cdxi7979m ^ cdxi7981m ^ cdxi5208m ^ cdxi5234m ^ cdxi7985m ^ cdxi5244m ^ cdxi7989m ^ cdxi5246m ^ cdxi8616m ^ cdxi5288m ^ cdxi5299m ^ cdxi8015m ^ cdxi5330m ^ cdxi5405m ^ cdxi9034m ^ cdxi5479m ^ cdxi8032m ^ cdxi5514m ^ cdxi8895m ^ cdxi5550m ^ cdxi5691m ^ cdxi5761m ^ cdxi5830m ^ cdxi5864m ^ cdxi5932m ^ cdxi5966m ^ cdxi5999m ^ cdxi8128m ^ cdxi6033m ^ cdxi8149m ^ cdxi8151m ^ cdxi9051m ^ cdxi8652m ^ cdxi6084m ^ cdxi8654m ^ cdxi8656m ^ cdxi8159m ^ cdxi6167m ^ cdxi6189m ^ cdxi8161m ^ cdxi6260m ^ cdxi6331m ^ cdxi8979m ^ cdxi6399m ^ cdxi6469m ^ cdxi6607m ^ cdxi6744m ^ cdxi8689m ^ cdxi7077m ^ cdxi7143m ^ cdxi7177m ^ cdxi8722m ^ cdxi7246m ^ cdxi7318m ^ cdxi7455m ^ cdxi9053m ^ r130m;
	reg_1_139 <= cdxi4663m ^ cdxi4678m ^ cdxi4683m ^ cdxi4688m ^ cdxi7789m ^ cdxi8554m ^ cdxi4694m ^ cdxi4697m ^ cdxi7791m ^ cdxi7793m ^ cdxi4703m ^ cdxi7797m ^ cdxi4707m ^ cdxi4709m ^ cdxi7799m ^ cdxi7801m ^ cdxi4736m ^ cdxi9013m ^ cdxi7822m ^ cdxi7830m ^ cdxi4747m ^ cdxi7835m ^ cdxi7837m ^ cdxi9015m ^ cdxi4756m ^ cdxi7843m ^ cdxi8563m ^ cdxi7849m ^ cdxi4811m ^ cdxi9017m ^ cdxi8572m ^ cdxi7853m ^ cdxi4829m ^ cdxi7855m ^ cdxi7857m ^ cdxi4848m ^ cdxi7859m ^ cdxi4853m ^ cdxi4859m ^ cdxi4861m ^ cdxi4865m ^ cdxi4867m ^ cdxi8862m ^ cdxi4871m ^ cdxi4883m ^ cdxi7886m ^ cdxi7902m ^ cdxi4943m ^ cdxi4962m ^ cdxi8585m ^ cdxi4999m ^ cdxi5017m ^ cdxi7927m ^ cdxi7936m ^ cdxi5036m ^ cdxi7961m ^ cdxi7979m ^ cdxi5162m ^ cdxi7981m ^ cdxi5179m ^ cdxi5217m ^ cdxi5234m ^ cdxi7985m ^ cdxi5244m ^ cdxi7987m ^ cdxi5246m ^ cdxi8614m ^ cdxi5248m ^ cdxi8616m ^ cdxi7991m ^ cdxi5267m ^ cdxi7993m ^ cdxi8002m ^ cdxi5288m ^ cdxi5299m ^ cdxi5309m ^ cdxi8015m ^ cdxi5330m ^ cdxi5367m ^ cdxi5442m ^ cdxi9034m ^ cdxi5479m ^ cdxi8032m ^ cdxi5514m ^ cdxi5550m ^ cdxi8927m ^ cdxi5586m ^ cdxi5657m ^ cdxi5691m ^ cdxi5761m ^ cdxi8064m ^ cdxi5830m ^ cdxi5864m ^ cdxi5932m ^ cdxi8096m ^ cdxi8145m ^ cdxi6033m ^ cdxi8147m ^ cdxi8153m ^ cdxi9051m ^ cdxi8652m ^ cdxi6084m ^ cdxi8155m ^ cdxi8656m ^ cdxi8157m ^ cdxi6185m ^ cdxi8161m ^ cdxi6206m ^ cdxi6331m ^ cdxi8979m ^ cdxi6399m ^ cdxi6537m ^ cdxi6607m ^ cdxi6676m ^ cdxi6812m ^ cdxi8689m ^ cdxi8258m ^ cdxi7177m ^ cdxi8722m ^ cdxi7246m ^ cdxi8724m ^ cdxi8357m ^ cdxi7455m ^ cdxi7722m ^ cdxi9053m ^ r131m;
	reg_1_140 <= cdxi9054m ^ cdxi4683m ^ cdxi7789m ^ cdxi4697m ^ cdxi7793m ^ cdxi8556m ^ cdxi7795m ^ cdxi7797m ^ cdxi4707m ^ cdxi4709m ^ cdxi7801m ^ cdxi4726m ^ cdxi9058m ^ cdxi4736m ^ cdxi4747m ^ cdxi7835m ^ cdxi9015m ^ cdxi4766m ^ cdxi7843m ^ cdxi4784m ^ cdxi7845m ^ cdxi8563m ^ cdxi7849m ^ cdxi4793m ^ cdxi4802m ^ cdxi8570m ^ cdxi8858m ^ cdxi9017m ^ cdxi7853m ^ cdxi4829m ^ cdxi4837m ^ cdxi4853m ^ cdxi4861m ^ cdxi8862m ^ cdxi4869m ^ cdxi4871m ^ cdxi4883m ^ cdxi7886m ^ cdxi4924m ^ cdxi7902m ^ cdxi7918m ^ cdxi8585m ^ cdxi4999m ^ cdxi8601m ^ cdxi5017m ^ cdxi7936m ^ cdxi5073m ^ cdxi7952m ^ cdxi5091m ^ cdxi7961m ^ cdxi5126m ^ cdxi5206m ^ cdxi5208m ^ cdxi5234m ^ cdxi7985m ^ cdxi7987m ^ cdxi5246m ^ cdxi5257m ^ cdxi8002m ^ cdxi5309m ^ cdxi8013m ^ cdxi8015m ^ cdxi5330m ^ cdxi5367m ^ cdxi5405m ^ cdxi5442m ^ cdxi5479m ^ cdxi8032m ^ cdxi5514m ^ cdxi8895m ^ cdxi5550m ^ cdxi8927m ^ cdxi5657m ^ cdxi8633m ^ cdxi5727m ^ cdxi5796m ^ cdxi5830m ^ cdxi5864m ^ cdxi5899m ^ cdxi5932m ^ cdxi5966m ^ cdxi5999m ^ cdxi8096m ^ cdxi8946m ^ cdxi6033m ^ cdxi8147m ^ cdxi8149m ^ cdxi8151m ^ cdxi9051m ^ cdxi6084m ^ cdxi8654m ^ cdxi8155m ^ cdxi8656m ^ cdxi6101m ^ cdxi8157m ^ cdxi6185m ^ cdxi6187m ^ cdxi6331m ^ cdxi8194m ^ cdxi6537m ^ cdxi6945m ^ cdxi7012m ^ cdxi7077m ^ cdxi7212m ^ cdxi8724m ^ cdxi8357m ^ cdxi9053m ^ cdxi8855m ^ r132m;
	reg_1_141 <= cdxi9063m ^ cdxi4663m ^ cdxi4683m ^ cdxi7789m ^ cdxi4694m ^ cdxi7791m ^ cdxi7793m ^ cdxi7795m ^ cdxi4707m ^ cdxi4709m ^ cdxi7806m ^ cdxi4716m ^ cdxi7814m ^ cdxi4736m ^ cdxi9013m ^ cdxi7822m ^ cdxi7835m ^ cdxi7839m ^ cdxi9015m ^ cdxi4756m ^ cdxi4766m ^ cdxi8563m ^ cdxi4802m ^ cdxi8570m ^ cdxi4811m ^ cdxi4820m ^ cdxi7851m ^ cdxi9017m ^ cdxi8574m ^ cdxi4829m ^ cdxi4835m ^ cdxi7857m ^ cdxi4837m ^ cdxi4848m ^ cdxi4853m ^ cdxi4861m ^ cdxi4863m ^ cdxi4867m ^ cdxi4871m ^ cdxi7861m ^ cdxi4883m ^ cdxi7918m ^ cdxi4943m ^ cdxi4981m ^ cdxi8585m ^ cdxi8601m ^ cdxi7927m ^ cdxi7952m ^ cdxi5091m ^ cdxi5109m ^ cdxi5144m ^ cdxi7979m ^ cdxi9064m ^ cdxi5162m ^ cdxi7981m ^ cdxi5208m ^ cdxi5234m ^ cdxi7985m ^ cdxi5244m ^ cdxi7987m ^ cdxi8614m ^ cdxi5248m ^ cdxi7993m ^ cdxi9066m ^ cdxi5288m ^ cdxi8013m ^ cdxi8015m ^ cdxi5330m ^ cdxi5442m ^ cdxi9034m ^ cdxi5479m ^ cdxi8032m ^ cdxi5514m ^ cdxi8895m ^ cdxi8927m ^ cdxi5657m ^ cdxi8633m ^ cdxi5796m ^ cdxi8944m ^ cdxi5899m ^ cdxi5932m ^ cdxi5966m ^ cdxi8096m ^ cdxi8128m ^ cdxi8650m ^ cdxi8149m ^ cdxi6066m ^ cdxi9068m ^ cdxi8153m ^ cdxi9051m ^ cdxi8652m ^ cdxi6084m ^ cdxi8155m ^ cdxi8656m ^ cdxi8157m ^ cdxi8159m ^ cdxi6167m ^ cdxi6189m ^ cdxi6206m ^ cdxi6260m ^ cdxi6399m ^ cdxi6469m ^ cdxi6676m ^ cdxi6744m ^ cdxi8258m ^ cdxi6945m ^ cdxi7077m ^ cdxi7143m ^ cdxi7177m ^ cdxi7246m ^ cdxi8724m ^ cdxi8357m ^ cdxi7455m ^ cdxi9053m ^ r133m;
end

assign x0 = cdxi132m ^ cdxi138m ^ cdxi144m ^ cdxi150m ^ cdxi156m ^ cdxi162m ^ cdxi164m ^ cdxi166m ^ cdxi172m ^ cdxi174m ^ cdxi176m ^ cdxi178m ^ cdxi180m ^ cdxi182m ^ cdxi194m ^ cdxi205m ^ cdxi216m ^ cdxi228m ^ cdxi238m ^ cdxi249m ^ cdxi259m ^ cdxi269m ^ cdxi279m ^ cdxi289m ^ cdxi299m ^ cdxi309m ^ cdxi319m ^ cdxi321m ^ cdxi323m ^ cdxi333m ^ cdxi335m ^ cdxi345m ^ cdxi347m ^ cdxi349m ^ cdxi351m ^ cdxi353m ^ cdxi355m ^ cdxi357m ^ cdxi359m ^ cdxi382m ^ cdxi403m ^ cdxi423m ^ cdxi443m ^ cdxi464m ^ cdxi483m ^ cdxi502m ^ cdxi522m ^ cdxi542m ^ cdxi560m ^ cdxi580m ^ cdxi599m ^ cdxi618m ^ cdxi636m ^ cdxi655m ^ cdxi674m ^ cdxi692m ^ cdxi710m ^ cdxi712m ^ cdxi714m ^ cdxi732m ^ cdxi750m ^ cdxi752m ^ cdxi754m ^ cdxi756m ^ cdxi774m ^ cdxi776m ^ cdxi794m ^ cdxi796m ^ cdxi798m ^ cdxi800m ^ cdxi818m ^ cdxi820m ^ cdxi859m ^ cdxi898m ^ cdxi936m ^ cdxi975m ^ cdxi1011m ^ cdxi1048m ^ cdxi1086m ^ cdxi1121m ^ cdxi1158m ^ cdxi1194m ^ cdxi1230m ^ cdxi1266m ^ cdxi1301m ^ cdxi1337m ^ cdxi1372m ^ cdxi1408m ^ cdxi1443m ^ cdxi1477m ^ cdxi1512m ^ cdxi1546m ^ cdxi1581m ^ cdxi1615m ^ cdxi1617m ^ cdxi1651m ^ cdxi1685m ^ cdxi1719m ^ cdxi1721m ^ cdxi1723m ^ cdxi1725m ^ cdxi1759m ^ cdxi1832m ^ cdxi1902m ^ cdxi1972m ^ cdxi2043m ^ cdxi2112m ^ cdxi2184m ^ cdxi2254m ^ cdxi2321m ^ cdxi2390m ^ cdxi2457m ^ cdxi2525m ^ cdxi2593m ^ cdxi2659m ^ cdxi2726m ^ cdxi2728m ^ cdxi2730m ^ cdxi2796m ^ cdxi2798m ^ cdxi2938m ^ cdxi3074m ^ cdxi3209m ^ cdxi3342m ^ reg_0_134;
assign y0 = cdxi144m ^ cdxi150m ^ cdxi156m ^ cdxi3345m ^ cdxi164m ^ cdxi172m ^ cdxi3347m ^ cdxi3349m ^ cdxi3351m ^ cdxi3353m ^ cdxi180m ^ cdxi3355m ^ cdxi3357m ^ cdxi3366m ^ cdxi205m ^ cdxi3375m ^ cdxi216m ^ cdxi3384m ^ cdxi3393m ^ cdxi228m ^ cdxi3395m ^ cdxi3397m ^ cdxi3399m ^ cdxi238m ^ cdxi249m ^ cdxi3401m ^ cdxi3403m ^ cdxi3405m ^ cdxi3407m ^ cdxi3409m ^ cdxi299m ^ cdxi3411m ^ cdxi3413m ^ cdxi319m ^ cdxi3415m ^ cdxi321m ^ cdxi3417m ^ cdxi3419m ^ cdxi347m ^ cdxi351m ^ cdxi353m ^ cdxi355m ^ cdxi357m ^ cdxi3421m ^ cdxi382m ^ cdxi3438m ^ cdxi403m ^ cdxi3455m ^ cdxi3472m ^ cdxi3489m ^ cdxi464m ^ cdxi483m ^ cdxi502m ^ cdxi522m ^ cdxi3491m ^ cdxi3508m ^ cdxi580m ^ cdxi3525m ^ cdxi618m ^ cdxi3527m ^ cdxi3544m ^ cdxi636m ^ cdxi3546m ^ cdxi3548m ^ cdxi692m ^ cdxi3550m ^ cdxi712m ^ cdxi750m ^ cdxi3552m ^ cdxi3554m ^ cdxi3556m ^ cdxi754m ^ cdxi774m ^ cdxi3558m ^ cdxi3560m ^ cdxi794m ^ cdxi3577m ^ cdxi3579m ^ cdxi798m ^ cdxi818m ^ cdxi3581m ^ cdxi3583m ^ cdxi859m ^ cdxi898m ^ cdxi1011m ^ cdxi3616m ^ cdxi1048m ^ cdxi1158m ^ cdxi1194m ^ cdxi1266m ^ cdxi3649m ^ cdxi1408m ^ cdxi3682m ^ cdxi3715m ^ cdxi3717m ^ cdxi3719m ^ cdxi3721m ^ cdxi3723m ^ cdxi3725m ^ cdxi1617m ^ cdxi3727m ^ cdxi1651m ^ cdxi3729m ^ cdxi3731m ^ cdxi1719m ^ cdxi1721m ^ cdxi1725m ^ cdxi3733m ^ cdxi1832m ^ cdxi1902m ^ cdxi1972m ^ cdxi2043m ^ cdxi3798m ^ cdxi2112m ^ cdxi2254m ^ cdxi2390m ^ cdxi2457m ^ cdxi3864m ^ cdxi2525m ^ cdxi2796m ^ cdxi2798m ^ cdxi3996m ^ cdxi3342m ^ cdxi4127m ^ reg_0_135;
assign z0 = cdxi132m ^ cdxi138m ^ cdxi144m ^ cdxi156m ^ cdxi164m ^ cdxi4130m ^ cdxi172m ^ cdxi4132m ^ cdxi4134m ^ cdxi178m ^ cdxi180m ^ cdxi182m ^ cdxi3366m ^ cdxi194m ^ cdxi216m ^ cdxi3393m ^ cdxi3395m ^ cdxi3397m ^ cdxi238m ^ cdxi3401m ^ cdxi3403m ^ cdxi269m ^ cdxi4143m ^ cdxi4145m ^ cdxi4147m ^ cdxi299m ^ cdxi3411m ^ cdxi4149m ^ cdxi4151m ^ cdxi3413m ^ cdxi319m ^ cdxi3417m ^ cdxi335m ^ cdxi3419m ^ cdxi345m ^ cdxi347m ^ cdxi349m ^ cdxi353m ^ cdxi4153m ^ cdxi3421m ^ cdxi382m ^ cdxi3472m ^ cdxi483m ^ cdxi4170m ^ cdxi502m ^ cdxi4187m ^ cdxi4189m ^ cdxi3491m ^ cdxi3508m ^ cdxi4191m ^ cdxi599m ^ cdxi618m ^ cdxi3544m ^ cdxi636m ^ cdxi655m ^ cdxi3546m ^ cdxi3548m ^ cdxi3550m ^ cdxi712m ^ cdxi732m ^ cdxi750m ^ cdxi3554m ^ cdxi754m ^ cdxi4193m ^ cdxi756m ^ cdxi4195m ^ cdxi3558m ^ cdxi3577m ^ cdxi800m ^ cdxi3581m ^ cdxi3583m ^ cdxi859m ^ cdxi936m ^ cdxi3616m ^ cdxi1086m ^ cdxi1121m ^ cdxi1158m ^ cdxi4228m ^ cdxi1266m ^ cdxi1301m ^ cdxi3649m ^ cdxi1337m ^ cdxi1443m ^ cdxi1546m ^ cdxi3715m ^ cdxi4230m ^ cdxi1581m ^ cdxi3721m ^ cdxi1615m ^ cdxi4232m ^ cdxi4234m ^ cdxi3727m ^ cdxi4236m ^ cdxi1685m ^ cdxi3731m ^ cdxi1721m ^ cdxi1723m ^ cdxi1725m ^ cdxi2043m ^ cdxi2184m ^ cdxi2254m ^ cdxi2321m ^ cdxi4301m ^ cdxi4303m ^ cdxi4305m ^ cdxi4435m ^ cdxi3209m ^ cdxi4127m ^ cdxi4437m ^ reg_0_136;
assign t0 = cdxi132m ^ cdxi138m ^ cdxi144m ^ cdxi156m ^ cdxi4130m ^ cdxi166m ^ cdxi172m ^ cdxi3347m ^ cdxi3349m ^ cdxi174m ^ cdxi176m ^ cdxi178m ^ cdxi182m ^ cdxi3355m ^ cdxi3357m ^ cdxi3366m ^ cdxi194m ^ cdxi205m ^ cdxi3375m ^ cdxi216m ^ cdxi3395m ^ cdxi238m ^ cdxi3401m ^ cdxi3403m ^ cdxi259m ^ cdxi4143m ^ cdxi3407m ^ cdxi4145m ^ cdxi279m ^ cdxi289m ^ cdxi4147m ^ cdxi299m ^ cdxi4440m ^ cdxi4442m ^ cdxi3413m ^ cdxi3415m ^ cdxi335m ^ cdxi349m ^ cdxi355m ^ cdxi4444m ^ cdxi359m ^ cdxi4461m ^ cdxi403m ^ cdxi3489m ^ cdxi4170m ^ cdxi522m ^ cdxi3491m ^ cdxi542m ^ cdxi560m ^ cdxi580m ^ cdxi4191m ^ cdxi3525m ^ cdxi636m ^ cdxi655m ^ cdxi674m ^ cdxi3548m ^ cdxi692m ^ cdxi3550m ^ cdxi714m ^ cdxi750m ^ cdxi4193m ^ cdxi756m ^ cdxi4195m ^ cdxi774m ^ cdxi3558m ^ cdxi3560m ^ cdxi798m ^ cdxi800m ^ cdxi820m ^ cdxi859m ^ cdxi898m ^ cdxi936m ^ cdxi975m ^ cdxi1011m ^ cdxi4494m ^ cdxi4527m ^ cdxi1121m ^ cdxi4529m ^ cdxi1372m ^ cdxi1408m ^ cdxi1443m ^ cdxi4531m ^ cdxi3719m ^ cdxi3721m ^ cdxi3723m ^ cdxi3725m ^ cdxi1617m ^ cdxi4236m ^ cdxi1651m ^ cdxi3731m ^ cdxi1719m ^ cdxi1721m ^ cdxi1725m ^ cdxi3733m ^ cdxi1759m ^ cdxi1832m ^ cdxi4596m ^ cdxi2043m ^ cdxi2112m ^ cdxi2184m ^ cdxi2254m ^ cdxi2321m ^ cdxi4301m ^ cdxi3864m ^ cdxi2525m ^ cdxi2659m ^ cdxi2726m ^ cdxi2728m ^ cdxi2796m ^ cdxi4303m ^ cdxi2798m ^ cdxi4305m ^ cdxi4435m ^ cdxi3209m ^ cdxi3342m ^ reg_0_137;
assign m0 = cdxi132m ^ cdxi138m ^ cdxi3345m ^ cdxi4130m ^ cdxi166m ^ cdxi172m ^ cdxi3349m ^ cdxi4132m ^ cdxi3351m ^ cdxi180m ^ cdxi182m ^ cdxi3366m ^ cdxi194m ^ cdxi205m ^ cdxi216m ^ cdxi4599m ^ cdxi3384m ^ cdxi228m ^ cdxi4601m ^ cdxi238m ^ cdxi249m ^ cdxi3401m ^ cdxi3405m ^ cdxi4143m ^ cdxi3407m ^ cdxi3409m ^ cdxi4145m ^ cdxi279m ^ cdxi289m ^ cdxi299m ^ cdxi4440m ^ cdxi4442m ^ cdxi3411m ^ cdxi4603m ^ cdxi4149m ^ cdxi4151m ^ cdxi3413m ^ cdxi319m ^ cdxi321m ^ cdxi3417m ^ cdxi335m ^ cdxi3419m ^ cdxi353m ^ cdxi355m ^ cdxi4444m ^ cdxi357m ^ cdxi4153m ^ cdxi3438m ^ cdxi4461m ^ cdxi3455m ^ cdxi423m ^ cdxi3472m ^ cdxi3508m ^ cdxi542m ^ cdxi560m ^ cdxi580m ^ cdxi3525m ^ cdxi599m ^ cdxi618m ^ cdxi3527m ^ cdxi655m ^ cdxi3546m ^ cdxi3548m ^ cdxi714m ^ cdxi750m ^ cdxi3552m ^ cdxi752m ^ cdxi3556m ^ cdxi754m ^ cdxi4195m ^ cdxi798m ^ cdxi818m ^ cdxi3583m ^ cdxi859m ^ cdxi936m ^ cdxi4636m ^ cdxi1011m ^ cdxi3616m ^ cdxi1048m ^ cdxi4494m ^ cdxi1086m ^ cdxi1230m ^ cdxi1301m ^ cdxi1372m ^ cdxi1408m ^ cdxi1477m ^ cdxi1512m ^ cdxi1546m ^ cdxi3715m ^ cdxi1581m ^ cdxi3721m ^ cdxi3723m ^ cdxi4638m ^ cdxi4232m ^ cdxi1617m ^ cdxi4234m ^ cdxi4236m ^ cdxi3731m ^ cdxi1719m ^ cdxi1725m ^ cdxi3733m ^ cdxi1832m ^ cdxi1902m ^ cdxi4596m ^ cdxi1972m ^ cdxi2043m ^ cdxi2184m ^ cdxi2321m ^ cdxi4301m ^ cdxi2659m ^ cdxi2726m ^ cdxi2728m ^ cdxi4303m ^ cdxi2798m ^ cdxi2938m ^ cdxi3074m ^ cdxi4127m ^ reg_0_138;
assign n0 = cdxi132m ^ cdxi150m ^ cdxi156m ^ cdxi162m ^ cdxi3345m ^ cdxi4130m ^ cdxi166m ^ cdxi172m ^ cdxi3347m ^ cdxi3349m ^ cdxi176m ^ cdxi3353m ^ cdxi180m ^ cdxi182m ^ cdxi3355m ^ cdxi3357m ^ cdxi216m ^ cdxi4599m ^ cdxi3384m ^ cdxi3393m ^ cdxi228m ^ cdxi3395m ^ cdxi3397m ^ cdxi4601m ^ cdxi238m ^ cdxi3403m ^ cdxi4143m ^ cdxi3409m ^ cdxi299m ^ cdxi4603m ^ cdxi4149m ^ cdxi3413m ^ cdxi319m ^ cdxi3415m ^ cdxi3417m ^ cdxi335m ^ cdxi3419m ^ cdxi345m ^ cdxi347m ^ cdxi349m ^ cdxi353m ^ cdxi355m ^ cdxi4444m ^ cdxi359m ^ cdxi382m ^ cdxi3455m ^ cdxi3472m ^ cdxi443m ^ cdxi464m ^ cdxi4170m ^ cdxi502m ^ cdxi522m ^ cdxi3491m ^ cdxi3508m ^ cdxi542m ^ cdxi3527m ^ cdxi3546m ^ cdxi674m ^ cdxi3548m ^ cdxi692m ^ cdxi732m ^ cdxi750m ^ cdxi3552m ^ cdxi752m ^ cdxi3554m ^ cdxi754m ^ cdxi4193m ^ cdxi756m ^ cdxi4195m ^ cdxi3558m ^ cdxi776m ^ cdxi3560m ^ cdxi3577m ^ cdxi798m ^ cdxi818m ^ cdxi820m ^ cdxi3583m ^ cdxi859m ^ cdxi898m ^ cdxi975m ^ cdxi4636m ^ cdxi1011m ^ cdxi3616m ^ cdxi1048m ^ cdxi1086m ^ cdxi4527m ^ cdxi1121m ^ cdxi1194m ^ cdxi1230m ^ cdxi1301m ^ cdxi3649m ^ cdxi1372m ^ cdxi1408m ^ cdxi1477m ^ cdxi3682m ^ cdxi3717m ^ cdxi1581m ^ cdxi3719m ^ cdxi3725m ^ cdxi4638m ^ cdxi4232m ^ cdxi1617m ^ cdxi3727m ^ cdxi4236m ^ cdxi3729m ^ cdxi1721m ^ cdxi3733m ^ cdxi1759m ^ cdxi1902m ^ cdxi4596m ^ cdxi1972m ^ cdxi2112m ^ cdxi2184m ^ cdxi2254m ^ cdxi2390m ^ cdxi4301m ^ cdxi3864m ^ cdxi2728m ^ cdxi4303m ^ cdxi2798m ^ cdxi4305m ^ cdxi3996m ^ cdxi3074m ^ cdxi3342m ^ cdxi4127m ^ reg_0_139;
assign p0 = cdxi156m ^ cdxi3345m ^ cdxi172m ^ cdxi3349m ^ cdxi4132m ^ cdxi3351m ^ cdxi3353m ^ cdxi180m ^ cdxi182m ^ cdxi3357m ^ cdxi205m ^ cdxi4649m ^ cdxi216m ^ cdxi228m ^ cdxi3395m ^ cdxi4601m ^ cdxi249m ^ cdxi3403m ^ cdxi269m ^ cdxi3405m ^ cdxi4143m ^ cdxi3409m ^ cdxi279m ^ cdxi289m ^ cdxi4147m ^ cdxi4440m ^ cdxi4603m ^ cdxi3413m ^ cdxi319m ^ cdxi323m ^ cdxi345m ^ cdxi349m ^ cdxi4444m ^ cdxi357m ^ cdxi359m ^ cdxi382m ^ cdxi3455m ^ cdxi423m ^ cdxi3472m ^ cdxi3489m ^ cdxi4170m ^ cdxi502m ^ cdxi4187m ^ cdxi522m ^ cdxi3508m ^ cdxi580m ^ cdxi3525m ^ cdxi599m ^ cdxi3527m ^ cdxi636m ^ cdxi712m ^ cdxi714m ^ cdxi750m ^ cdxi3552m ^ cdxi3554m ^ cdxi754m ^ cdxi774m ^ cdxi3577m ^ cdxi820m ^ cdxi3581m ^ cdxi3583m ^ cdxi859m ^ cdxi898m ^ cdxi936m ^ cdxi975m ^ cdxi1011m ^ cdxi3616m ^ cdxi1048m ^ cdxi4494m ^ cdxi1086m ^ cdxi4527m ^ cdxi1194m ^ cdxi4228m ^ cdxi1266m ^ cdxi1337m ^ cdxi1372m ^ cdxi1408m ^ cdxi1443m ^ cdxi1477m ^ cdxi1512m ^ cdxi1546m ^ cdxi3682m ^ cdxi4531m ^ cdxi1581m ^ cdxi3719m ^ cdxi3721m ^ cdxi3723m ^ cdxi4638m ^ cdxi1617m ^ cdxi4234m ^ cdxi3727m ^ cdxi4236m ^ cdxi1651m ^ cdxi3729m ^ cdxi1721m ^ cdxi1723m ^ cdxi1902m ^ cdxi3798m ^ cdxi2112m ^ cdxi2525m ^ cdxi2593m ^ cdxi2659m ^ cdxi2796m ^ cdxi4305m ^ cdxi3996m ^ cdxi4127m ^ cdxi4437m ^ reg_0_140;
assign q0 = cdxi132m ^ cdxi156m ^ cdxi3345m ^ cdxi166m ^ cdxi3347m ^ cdxi3349m ^ cdxi3351m ^ cdxi180m ^ cdxi182m ^ cdxi3366m ^ cdxi194m ^ cdxi3375m ^ cdxi216m ^ cdxi4599m ^ cdxi3384m ^ cdxi3395m ^ cdxi3399m ^ cdxi4601m ^ cdxi238m ^ cdxi249m ^ cdxi4143m ^ cdxi289m ^ cdxi4147m ^ cdxi299m ^ cdxi309m ^ cdxi3411m ^ cdxi4603m ^ cdxi4151m ^ cdxi319m ^ cdxi321m ^ cdxi3417m ^ cdxi323m ^ cdxi335m ^ cdxi345m ^ cdxi349m ^ cdxi351m ^ cdxi355m ^ cdxi359m ^ cdxi3421m ^ cdxi382m ^ cdxi3489m ^ cdxi443m ^ cdxi483m ^ cdxi4170m ^ cdxi4187m ^ cdxi3491m ^ cdxi3525m ^ cdxi599m ^ cdxi618m ^ cdxi655m ^ cdxi3546m ^ cdxi4652m ^ cdxi674m ^ cdxi3548m ^ cdxi714m ^ cdxi750m ^ cdxi3552m ^ cdxi752m ^ cdxi3554m ^ cdxi4193m ^ cdxi756m ^ cdxi3560m ^ cdxi4654m ^ cdxi798m ^ cdxi3581m ^ cdxi3583m ^ cdxi859m ^ cdxi975m ^ cdxi4636m ^ cdxi1011m ^ cdxi3616m ^ cdxi1048m ^ cdxi4494m ^ cdxi4527m ^ cdxi1194m ^ cdxi4228m ^ cdxi1337m ^ cdxi4529m ^ cdxi1443m ^ cdxi1477m ^ cdxi1512m ^ cdxi3682m ^ cdxi3715m ^ cdxi4230m ^ cdxi3721m ^ cdxi1615m ^ cdxi4656m ^ cdxi3725m ^ cdxi4638m ^ cdxi4232m ^ cdxi1617m ^ cdxi3727m ^ cdxi4236m ^ cdxi3729m ^ cdxi3731m ^ cdxi1719m ^ cdxi1725m ^ cdxi1759m ^ cdxi1832m ^ cdxi1972m ^ cdxi2043m ^ cdxi2254m ^ cdxi2321m ^ cdxi3864m ^ cdxi2525m ^ cdxi2659m ^ cdxi2726m ^ cdxi2728m ^ cdxi2798m ^ cdxi4305m ^ cdxi3996m ^ cdxi3074m ^ cdxi4127m ^ reg_0_141;



assign x1 = cdxi4666m ^ cdxi4671m ^ cdxi4676m ^ cdxi4681m ^ cdxi4686m ^ cdxi4691m ^ cdxi4693m ^ cdxi4695m ^ cdxi4700m ^ cdxi4702m ^ cdxi4704m ^ cdxi4706m ^ cdxi4708m ^ cdxi4710m ^ cdxi4721m ^ cdxi4731m ^ cdxi4741m ^ cdxi4752m ^ cdxi4761m ^ cdxi4771m ^ cdxi4780m ^ cdxi4789m ^ cdxi4798m ^ cdxi4807m ^ cdxi4816m ^ cdxi4825m ^ cdxi4834m ^ cdxi4836m ^ cdxi4838m ^ cdxi4847m ^ cdxi4849m ^ cdxi4858m ^ cdxi4860m ^ cdxi4862m ^ cdxi4864m ^ cdxi4866m ^ cdxi4868m ^ cdxi4870m ^ cdxi4872m ^ cdxi4894m ^ cdxi4914m ^ cdxi4933m ^ cdxi4952m ^ cdxi4972m ^ cdxi4990m ^ cdxi5008m ^ cdxi5027m ^ cdxi5046m ^ cdxi5063m ^ cdxi5082m ^ cdxi5100m ^ cdxi5118m ^ cdxi5135m ^ cdxi5153m ^ cdxi5171m ^ cdxi5188m ^ cdxi5205m ^ cdxi5207m ^ cdxi5209m ^ cdxi5226m ^ cdxi5243m ^ cdxi5245m ^ cdxi5247m ^ cdxi5249m ^ cdxi5266m ^ cdxi5268m ^ cdxi5285m ^ cdxi5287m ^ cdxi5289m ^ cdxi5291m ^ cdxi5308m ^ cdxi5310m ^ cdxi5348m ^ cdxi5386m ^ cdxi5423m ^ cdxi5461m ^ cdxi5496m ^ cdxi5532m ^ cdxi5569m ^ cdxi5603m ^ cdxi5639m ^ cdxi5674m ^ cdxi5709m ^ cdxi5744m ^ cdxi5778m ^ cdxi5813m ^ cdxi5847m ^ cdxi5882m ^ cdxi5916m ^ cdxi5949m ^ cdxi5983m ^ cdxi6016m ^ cdxi6050m ^ cdxi6083m ^ cdxi6085m ^ cdxi6118m ^ cdxi6151m ^ cdxi6184m ^ cdxi6186m ^ cdxi6188m ^ cdxi6190m ^ cdxi6223m ^ cdxi6295m ^ cdxi6364m ^ cdxi6433m ^ cdxi6503m ^ cdxi6571m ^ cdxi6642m ^ cdxi6711m ^ cdxi6777m ^ cdxi6845m ^ cdxi6911m ^ cdxi6978m ^ cdxi7045m ^ cdxi7110m ^ cdxi7176m ^ cdxi7178m ^ cdxi7180m ^ cdxi7245m ^ cdxi7247m ^ cdxi7386m ^ cdxi7521m ^ cdxi7655m ^ cdxi7787m ^ reg_1_134;
assign y1 = cdxi4676m ^ cdxi4681m ^ cdxi4686m ^ cdxi7790m ^ cdxi4693m ^ cdxi4700m ^ cdxi7792m ^ cdxi7794m ^ cdxi7796m ^ cdxi7798m ^ cdxi4708m ^ cdxi7800m ^ cdxi7802m ^ cdxi7810m ^ cdxi4731m ^ cdxi7818m ^ cdxi4741m ^ cdxi7826m ^ cdxi7834m ^ cdxi4752m ^ cdxi7836m ^ cdxi7838m ^ cdxi7840m ^ cdxi4761m ^ cdxi4771m ^ cdxi7842m ^ cdxi7844m ^ cdxi7846m ^ cdxi7848m ^ cdxi7850m ^ cdxi4816m ^ cdxi7852m ^ cdxi7854m ^ cdxi4834m ^ cdxi7856m ^ cdxi4836m ^ cdxi7858m ^ cdxi7860m ^ cdxi4860m ^ cdxi4864m ^ cdxi4866m ^ cdxi4868m ^ cdxi4870m ^ cdxi7862m ^ cdxi4894m ^ cdxi7878m ^ cdxi4914m ^ cdxi7894m ^ cdxi7910m ^ cdxi7926m ^ cdxi4972m ^ cdxi4990m ^ cdxi5008m ^ cdxi5027m ^ cdxi7928m ^ cdxi7944m ^ cdxi5082m ^ cdxi7960m ^ cdxi5118m ^ cdxi7962m ^ cdxi7978m ^ cdxi5135m ^ cdxi7980m ^ cdxi7982m ^ cdxi5188m ^ cdxi7984m ^ cdxi5207m ^ cdxi5243m ^ cdxi7986m ^ cdxi7988m ^ cdxi7990m ^ cdxi5247m ^ cdxi5266m ^ cdxi7992m ^ cdxi7994m ^ cdxi5285m ^ cdxi8010m ^ cdxi8012m ^ cdxi5289m ^ cdxi5308m ^ cdxi8014m ^ cdxi8016m ^ cdxi5348m ^ cdxi5386m ^ cdxi5496m ^ cdxi8048m ^ cdxi5532m ^ cdxi5639m ^ cdxi5674m ^ cdxi5744m ^ cdxi8080m ^ cdxi5882m ^ cdxi8112m ^ cdxi8144m ^ cdxi8146m ^ cdxi8148m ^ cdxi8150m ^ cdxi8152m ^ cdxi8154m ^ cdxi6085m ^ cdxi8156m ^ cdxi6118m ^ cdxi8158m ^ cdxi8160m ^ cdxi6184m ^ cdxi6186m ^ cdxi6190m ^ cdxi8162m ^ cdxi6295m ^ cdxi6364m ^ cdxi6433m ^ cdxi6503m ^ cdxi8226m ^ cdxi6571m ^ cdxi6711m ^ cdxi6845m ^ cdxi6911m ^ cdxi8291m ^ cdxi6978m ^ cdxi7245m ^ cdxi7247m ^ cdxi8422m ^ cdxi7787m ^ cdxi8552m ^ reg_1_135;
assign z1 = cdxi4666m ^ cdxi4671m ^ cdxi4676m ^ cdxi4686m ^ cdxi4693m ^ cdxi8555m ^ cdxi4700m ^ cdxi8557m ^ cdxi8559m ^ cdxi4706m ^ cdxi4708m ^ cdxi4710m ^ cdxi7810m ^ cdxi4721m ^ cdxi4741m ^ cdxi7834m ^ cdxi7836m ^ cdxi7838m ^ cdxi4761m ^ cdxi7842m ^ cdxi7844m ^ cdxi4789m ^ cdxi8567m ^ cdxi8569m ^ cdxi8571m ^ cdxi4816m ^ cdxi7852m ^ cdxi8573m ^ cdxi8575m ^ cdxi7854m ^ cdxi4834m ^ cdxi7858m ^ cdxi4849m ^ cdxi7860m ^ cdxi4858m ^ cdxi4860m ^ cdxi4862m ^ cdxi4866m ^ cdxi8577m ^ cdxi7862m ^ cdxi4894m ^ cdxi7910m ^ cdxi4990m ^ cdxi8593m ^ cdxi5008m ^ cdxi8609m ^ cdxi8611m ^ cdxi7928m ^ cdxi7944m ^ cdxi8613m ^ cdxi5100m ^ cdxi5118m ^ cdxi7978m ^ cdxi5135m ^ cdxi5153m ^ cdxi7980m ^ cdxi7982m ^ cdxi7984m ^ cdxi5207m ^ cdxi5226m ^ cdxi5243m ^ cdxi7988m ^ cdxi5247m ^ cdxi8615m ^ cdxi5249m ^ cdxi8617m ^ cdxi7992m ^ cdxi8010m ^ cdxi5291m ^ cdxi8014m ^ cdxi8016m ^ cdxi5348m ^ cdxi5423m ^ cdxi8048m ^ cdxi5569m ^ cdxi5603m ^ cdxi5639m ^ cdxi8649m ^ cdxi5744m ^ cdxi5778m ^ cdxi8080m ^ cdxi5813m ^ cdxi5916m ^ cdxi6016m ^ cdxi8144m ^ cdxi8651m ^ cdxi6050m ^ cdxi8150m ^ cdxi6083m ^ cdxi8653m ^ cdxi8655m ^ cdxi8156m ^ cdxi8657m ^ cdxi6151m ^ cdxi8160m ^ cdxi6186m ^ cdxi6188m ^ cdxi6190m ^ cdxi6503m ^ cdxi6642m ^ cdxi6711m ^ cdxi6777m ^ cdxi8721m ^ cdxi8723m ^ cdxi8725m ^ cdxi8854m ^ cdxi7655m ^ cdxi8552m ^ cdxi8856m ^ reg_1_136;
assign t1 = cdxi4666m ^ cdxi4671m ^ cdxi4676m ^ cdxi4686m ^ cdxi8555m ^ cdxi4695m ^ cdxi4700m ^ cdxi7792m ^ cdxi7794m ^ cdxi4702m ^ cdxi4704m ^ cdxi4706m ^ cdxi4710m ^ cdxi7800m ^ cdxi7802m ^ cdxi7810m ^ cdxi4721m ^ cdxi4731m ^ cdxi7818m ^ cdxi4741m ^ cdxi7836m ^ cdxi4761m ^ cdxi7842m ^ cdxi7844m ^ cdxi4780m ^ cdxi8567m ^ cdxi7848m ^ cdxi8569m ^ cdxi4798m ^ cdxi4807m ^ cdxi8571m ^ cdxi4816m ^ cdxi8859m ^ cdxi8861m ^ cdxi7854m ^ cdxi7856m ^ cdxi4849m ^ cdxi4862m ^ cdxi4868m ^ cdxi8863m ^ cdxi4872m ^ cdxi8879m ^ cdxi4914m ^ cdxi7926m ^ cdxi8593m ^ cdxi5027m ^ cdxi7928m ^ cdxi5046m ^ cdxi5063m ^ cdxi5082m ^ cdxi8613m ^ cdxi7960m ^ cdxi5135m ^ cdxi5153m ^ cdxi5171m ^ cdxi7982m ^ cdxi5188m ^ cdxi7984m ^ cdxi5209m ^ cdxi5243m ^ cdxi8615m ^ cdxi5249m ^ cdxi8617m ^ cdxi5266m ^ cdxi7992m ^ cdxi7994m ^ cdxi5289m ^ cdxi5291m ^ cdxi5310m ^ cdxi5348m ^ cdxi5386m ^ cdxi5423m ^ cdxi5461m ^ cdxi5496m ^ cdxi8911m ^ cdxi8943m ^ cdxi5603m ^ cdxi8945m ^ cdxi5847m ^ cdxi5882m ^ cdxi5916m ^ cdxi8947m ^ cdxi8148m ^ cdxi8150m ^ cdxi8152m ^ cdxi8154m ^ cdxi6085m ^ cdxi8657m ^ cdxi6118m ^ cdxi8160m ^ cdxi6184m ^ cdxi6186m ^ cdxi6190m ^ cdxi8162m ^ cdxi6223m ^ cdxi6295m ^ cdxi9011m ^ cdxi6503m ^ cdxi6571m ^ cdxi6642m ^ cdxi6711m ^ cdxi6777m ^ cdxi8721m ^ cdxi8291m ^ cdxi6978m ^ cdxi7110m ^ cdxi7176m ^ cdxi7178m ^ cdxi7245m ^ cdxi8723m ^ cdxi7247m ^ cdxi8725m ^ cdxi8854m ^ cdxi7655m ^ cdxi7787m ^ reg_1_137;
assign m1 = cdxi4666m ^ cdxi4671m ^ cdxi7790m ^ cdxi8555m ^ cdxi4695m ^ cdxi4700m ^ cdxi7794m ^ cdxi8557m ^ cdxi7796m ^ cdxi4708m ^ cdxi4710m ^ cdxi7810m ^ cdxi4721m ^ cdxi4731m ^ cdxi4741m ^ cdxi9014m ^ cdxi7826m ^ cdxi4752m ^ cdxi9016m ^ cdxi4761m ^ cdxi4771m ^ cdxi7842m ^ cdxi7846m ^ cdxi8567m ^ cdxi7848m ^ cdxi7850m ^ cdxi8569m ^ cdxi4798m ^ cdxi4807m ^ cdxi4816m ^ cdxi8859m ^ cdxi8861m ^ cdxi7852m ^ cdxi9018m ^ cdxi8573m ^ cdxi8575m ^ cdxi7854m ^ cdxi4834m ^ cdxi4836m ^ cdxi7858m ^ cdxi4849m ^ cdxi7860m ^ cdxi4866m ^ cdxi4868m ^ cdxi8863m ^ cdxi4870m ^ cdxi8577m ^ cdxi7878m ^ cdxi8879m ^ cdxi7894m ^ cdxi4933m ^ cdxi7910m ^ cdxi7944m ^ cdxi5046m ^ cdxi5063m ^ cdxi5082m ^ cdxi7960m ^ cdxi5100m ^ cdxi5118m ^ cdxi7962m ^ cdxi5153m ^ cdxi7980m ^ cdxi7982m ^ cdxi5209m ^ cdxi5243m ^ cdxi7986m ^ cdxi5245m ^ cdxi7990m ^ cdxi5247m ^ cdxi8617m ^ cdxi5289m ^ cdxi5308m ^ cdxi8016m ^ cdxi5348m ^ cdxi5423m ^ cdxi9050m ^ cdxi5496m ^ cdxi8048m ^ cdxi5532m ^ cdxi8911m ^ cdxi5569m ^ cdxi5709m ^ cdxi5778m ^ cdxi5847m ^ cdxi5882m ^ cdxi5949m ^ cdxi5983m ^ cdxi6016m ^ cdxi8144m ^ cdxi6050m ^ cdxi8150m ^ cdxi8152m ^ cdxi9052m ^ cdxi8653m ^ cdxi6085m ^ cdxi8655m ^ cdxi8657m ^ cdxi8160m ^ cdxi6184m ^ cdxi6190m ^ cdxi8162m ^ cdxi6295m ^ cdxi6364m ^ cdxi9011m ^ cdxi6433m ^ cdxi6503m ^ cdxi6642m ^ cdxi6777m ^ cdxi8721m ^ cdxi7110m ^ cdxi7176m ^ cdxi7178m ^ cdxi8723m ^ cdxi7247m ^ cdxi7386m ^ cdxi7521m ^ cdxi8552m ^ reg_1_138;
assign n1 = cdxi4666m ^ cdxi4681m ^ cdxi4686m ^ cdxi4691m ^ cdxi7790m ^ cdxi8555m ^ cdxi4695m ^ cdxi4700m ^ cdxi7792m ^ cdxi7794m ^ cdxi4704m ^ cdxi7798m ^ cdxi4708m ^ cdxi4710m ^ cdxi7800m ^ cdxi7802m ^ cdxi4741m ^ cdxi9014m ^ cdxi7826m ^ cdxi7834m ^ cdxi4752m ^ cdxi7836m ^ cdxi7838m ^ cdxi9016m ^ cdxi4761m ^ cdxi7844m ^ cdxi8567m ^ cdxi7850m ^ cdxi4816m ^ cdxi9018m ^ cdxi8573m ^ cdxi7854m ^ cdxi4834m ^ cdxi7856m ^ cdxi7858m ^ cdxi4849m ^ cdxi7860m ^ cdxi4858m ^ cdxi4860m ^ cdxi4862m ^ cdxi4866m ^ cdxi4868m ^ cdxi8863m ^ cdxi4872m ^ cdxi4894m ^ cdxi7894m ^ cdxi7910m ^ cdxi4952m ^ cdxi4972m ^ cdxi8593m ^ cdxi5008m ^ cdxi5027m ^ cdxi7928m ^ cdxi7944m ^ cdxi5046m ^ cdxi7962m ^ cdxi7980m ^ cdxi5171m ^ cdxi7982m ^ cdxi5188m ^ cdxi5226m ^ cdxi5243m ^ cdxi7986m ^ cdxi5245m ^ cdxi7988m ^ cdxi5247m ^ cdxi8615m ^ cdxi5249m ^ cdxi8617m ^ cdxi7992m ^ cdxi5268m ^ cdxi7994m ^ cdxi8010m ^ cdxi5289m ^ cdxi5308m ^ cdxi5310m ^ cdxi8016m ^ cdxi5348m ^ cdxi5386m ^ cdxi5461m ^ cdxi9050m ^ cdxi5496m ^ cdxi8048m ^ cdxi5532m ^ cdxi5569m ^ cdxi8943m ^ cdxi5603m ^ cdxi5674m ^ cdxi5709m ^ cdxi5778m ^ cdxi8080m ^ cdxi5847m ^ cdxi5882m ^ cdxi5949m ^ cdxi8112m ^ cdxi8146m ^ cdxi6050m ^ cdxi8148m ^ cdxi8154m ^ cdxi9052m ^ cdxi8653m ^ cdxi6085m ^ cdxi8156m ^ cdxi8657m ^ cdxi8158m ^ cdxi6186m ^ cdxi8162m ^ cdxi6223m ^ cdxi6364m ^ cdxi9011m ^ cdxi6433m ^ cdxi6571m ^ cdxi6642m ^ cdxi6711m ^ cdxi6845m ^ cdxi8721m ^ cdxi8291m ^ cdxi7178m ^ cdxi8723m ^ cdxi7247m ^ cdxi8725m ^ cdxi8422m ^ cdxi7521m ^ cdxi7787m ^ cdxi8552m ^ reg_1_139;
assign p1 = cdxi4686m ^ cdxi7790m ^ cdxi4700m ^ cdxi7794m ^ cdxi8557m ^ cdxi7796m ^ cdxi7798m ^ cdxi4708m ^ cdxi4710m ^ cdxi7802m ^ cdxi4731m ^ cdxi9062m ^ cdxi4741m ^ cdxi4752m ^ cdxi7836m ^ cdxi9016m ^ cdxi4771m ^ cdxi7844m ^ cdxi4789m ^ cdxi7846m ^ cdxi8567m ^ cdxi7850m ^ cdxi4798m ^ cdxi4807m ^ cdxi8571m ^ cdxi8859m ^ cdxi9018m ^ cdxi7854m ^ cdxi4834m ^ cdxi4838m ^ cdxi4858m ^ cdxi4862m ^ cdxi8863m ^ cdxi4870m ^ cdxi4872m ^ cdxi4894m ^ cdxi7894m ^ cdxi4933m ^ cdxi7910m ^ cdxi7926m ^ cdxi8593m ^ cdxi5008m ^ cdxi8609m ^ cdxi5027m ^ cdxi7944m ^ cdxi5082m ^ cdxi7960m ^ cdxi5100m ^ cdxi7962m ^ cdxi5135m ^ cdxi5207m ^ cdxi5209m ^ cdxi5243m ^ cdxi7986m ^ cdxi7988m ^ cdxi5247m ^ cdxi5266m ^ cdxi8010m ^ cdxi5310m ^ cdxi8014m ^ cdxi8016m ^ cdxi5348m ^ cdxi5386m ^ cdxi5423m ^ cdxi5461m ^ cdxi5496m ^ cdxi8048m ^ cdxi5532m ^ cdxi8911m ^ cdxi5569m ^ cdxi8943m ^ cdxi5674m ^ cdxi8649m ^ cdxi5744m ^ cdxi5813m ^ cdxi5847m ^ cdxi5882m ^ cdxi5916m ^ cdxi5949m ^ cdxi5983m ^ cdxi6016m ^ cdxi8112m ^ cdxi8947m ^ cdxi6050m ^ cdxi8148m ^ cdxi8150m ^ cdxi8152m ^ cdxi9052m ^ cdxi6085m ^ cdxi8655m ^ cdxi8156m ^ cdxi8657m ^ cdxi6118m ^ cdxi8158m ^ cdxi6186m ^ cdxi6188m ^ cdxi6364m ^ cdxi8226m ^ cdxi6571m ^ cdxi6978m ^ cdxi7045m ^ cdxi7110m ^ cdxi7245m ^ cdxi8725m ^ cdxi8422m ^ cdxi8552m ^ cdxi8856m ^ reg_1_140;
assign q1 = cdxi4666m ^ cdxi4686m ^ cdxi7790m ^ cdxi4695m ^ cdxi7792m ^ cdxi7794m ^ cdxi7796m ^ cdxi4708m ^ cdxi4710m ^ cdxi7810m ^ cdxi4721m ^ cdxi7818m ^ cdxi4741m ^ cdxi9014m ^ cdxi7826m ^ cdxi7836m ^ cdxi7840m ^ cdxi9016m ^ cdxi4761m ^ cdxi4771m ^ cdxi8567m ^ cdxi4807m ^ cdxi8571m ^ cdxi4816m ^ cdxi4825m ^ cdxi7852m ^ cdxi9018m ^ cdxi8575m ^ cdxi4834m ^ cdxi4836m ^ cdxi7858m ^ cdxi4838m ^ cdxi4849m ^ cdxi4858m ^ cdxi4862m ^ cdxi4864m ^ cdxi4868m ^ cdxi4872m ^ cdxi7862m ^ cdxi4894m ^ cdxi7926m ^ cdxi4952m ^ cdxi4990m ^ cdxi8593m ^ cdxi8609m ^ cdxi7928m ^ cdxi7960m ^ cdxi5100m ^ cdxi5118m ^ cdxi5153m ^ cdxi7980m ^ cdxi9065m ^ cdxi5171m ^ cdxi7982m ^ cdxi5209m ^ cdxi5243m ^ cdxi7986m ^ cdxi5245m ^ cdxi7988m ^ cdxi8615m ^ cdxi5249m ^ cdxi7994m ^ cdxi9067m ^ cdxi5289m ^ cdxi8014m ^ cdxi8016m ^ cdxi5348m ^ cdxi5461m ^ cdxi9050m ^ cdxi5496m ^ cdxi8048m ^ cdxi5532m ^ cdxi8911m ^ cdxi8943m ^ cdxi5674m ^ cdxi8649m ^ cdxi5813m ^ cdxi8945m ^ cdxi5916m ^ cdxi5949m ^ cdxi5983m ^ cdxi8112m ^ cdxi8144m ^ cdxi8651m ^ cdxi8150m ^ cdxi6083m ^ cdxi9069m ^ cdxi8154m ^ cdxi9052m ^ cdxi8653m ^ cdxi6085m ^ cdxi8156m ^ cdxi8657m ^ cdxi8158m ^ cdxi8160m ^ cdxi6184m ^ cdxi6190m ^ cdxi6223m ^ cdxi6295m ^ cdxi6433m ^ cdxi6503m ^ cdxi6711m ^ cdxi6777m ^ cdxi8291m ^ cdxi6978m ^ cdxi7110m ^ cdxi7176m ^ cdxi7178m ^ cdxi7247m ^ cdxi8725m ^ cdxi8422m ^ cdxi7521m ^ cdxi8552m ^ reg_1_141;



assign x0y0z0t0m0n0p0q0 = {q0,p0,n0,m0,t0,z0,y0,x0};
assign x1y1z1t1m1n1p1q1 = {q1,p1,n1,m1,t1,z1,y1,x1};

wire [7:0] AT2in0, AT2in1, AT2out0, AT2out1;

assign AT2in0 = x0y0z0t0m0n0p0q0;
assign AT2in1 = x1y1z1t1m1n1p1q1;



wire [7:0] matrix1[0:7];
assign {matrix1[0], matrix1[1], matrix1[2], matrix1[3], matrix1[4], matrix1[5], matrix1[6], matrix1[7]} = { 8'h88 ,8'hA9 ,8'h4B ,8'h11 ,8'h68 ,8'h5D ,8'h83 ,8'h3F };
wire [7:0] constant1 = 8'h21 ;

assign AT2out0[7:7] = (matrix1[0][7:7]&AT2in0[7:7]) ^ (matrix1[0][6:6]&AT2in0[6:6]) ^ (matrix1[0][5:5]&AT2in0[5:5]) ^ (matrix1[0][4:4]&AT2in0[4:4]) ^ (matrix1[0][3:3]&AT2in0[3:3]) ^ (matrix1[0][2:2]&AT2in0[2:2]) ^ (matrix1[0][1:1]&AT2in0[1:1]) ^ (matrix1[0][0:0]&AT2in0[0:0]) ^ constant1[7:7]; 
assign AT2out0[6:6] = (matrix1[1][7:7]&AT2in0[7:7]) ^ (matrix1[1][6:6]&AT2in0[6:6]) ^ (matrix1[1][5:5]&AT2in0[5:5]) ^ (matrix1[1][4:4]&AT2in0[4:4]) ^ (matrix1[1][3:3]&AT2in0[3:3]) ^ (matrix1[1][2:2]&AT2in0[2:2]) ^ (matrix1[1][1:1]&AT2in0[1:1]) ^ (matrix1[1][0:0]&AT2in0[0:0]) ^ constant1[6:6]; 
assign AT2out0[5:5] = (matrix1[2][7:7]&AT2in0[7:7]) ^ (matrix1[2][6:6]&AT2in0[6:6]) ^ (matrix1[2][5:5]&AT2in0[5:5]) ^ (matrix1[2][4:4]&AT2in0[4:4]) ^ (matrix1[2][3:3]&AT2in0[3:3]) ^ (matrix1[2][2:2]&AT2in0[2:2]) ^ (matrix1[2][1:1]&AT2in0[1:1]) ^ (matrix1[2][0:0]&AT2in0[0:0]) ^ constant1[5:5]; 
assign AT2out0[4:4] = (matrix1[3][7:7]&AT2in0[7:7]) ^ (matrix1[3][6:6]&AT2in0[6:6]) ^ (matrix1[3][5:5]&AT2in0[5:5]) ^ (matrix1[3][4:4]&AT2in0[4:4]) ^ (matrix1[3][3:3]&AT2in0[3:3]) ^ (matrix1[3][2:2]&AT2in0[2:2]) ^ (matrix1[3][1:1]&AT2in0[1:1]) ^ (matrix1[3][0:0]&AT2in0[0:0]) ^ constant1[4:4]; 
assign AT2out0[3:3] = (matrix1[4][7:7]&AT2in0[7:7]) ^ (matrix1[4][6:6]&AT2in0[6:6]) ^ (matrix1[4][5:5]&AT2in0[5:5]) ^ (matrix1[4][4:4]&AT2in0[4:4]) ^ (matrix1[4][3:3]&AT2in0[3:3]) ^ (matrix1[4][2:2]&AT2in0[2:2]) ^ (matrix1[4][1:1]&AT2in0[1:1]) ^ (matrix1[4][0:0]&AT2in0[0:0]) ^ constant1[3:3]; 
assign AT2out0[2:2] = (matrix1[5][7:7]&AT2in0[7:7]) ^ (matrix1[5][6:6]&AT2in0[6:6]) ^ (matrix1[5][5:5]&AT2in0[5:5]) ^ (matrix1[5][4:4]&AT2in0[4:4]) ^ (matrix1[5][3:3]&AT2in0[3:3]) ^ (matrix1[5][2:2]&AT2in0[2:2]) ^ (matrix1[5][1:1]&AT2in0[1:1]) ^ (matrix1[5][0:0]&AT2in0[0:0]) ^ constant1[2:2]; 
assign AT2out0[1:1] = (matrix1[6][7:7]&AT2in0[7:7]) ^ (matrix1[6][6:6]&AT2in0[6:6]) ^ (matrix1[6][5:5]&AT2in0[5:5]) ^ (matrix1[6][4:4]&AT2in0[4:4]) ^ (matrix1[6][3:3]&AT2in0[3:3]) ^ (matrix1[6][2:2]&AT2in0[2:2]) ^ (matrix1[6][1:1]&AT2in0[1:1]) ^ (matrix1[6][0:0]&AT2in0[0:0]) ^ constant1[1:1]; 
assign AT2out0[0:0] = (matrix1[7][7:7]&AT2in0[7:7]) ^ (matrix1[7][6:6]&AT2in0[6:6]) ^ (matrix1[7][5:5]&AT2in0[5:5]) ^ (matrix1[7][4:4]&AT2in0[4:4]) ^ (matrix1[7][3:3]&AT2in0[3:3]) ^ (matrix1[7][2:2]&AT2in0[2:2]) ^ (matrix1[7][1:1]&AT2in0[1:1]) ^ (matrix1[7][0:0]&AT2in0[0:0]) ^ constant1[0:0]; 


assign AT2out1[7:7] = (matrix1[0][7:7]&AT2in1[7:7]) ^ (matrix1[0][6:6]&AT2in1[6:6]) ^ (matrix1[0][5:5]&AT2in1[5:5]) ^ (matrix1[0][4:4]&AT2in1[4:4]) ^ (matrix1[0][3:3]&AT2in1[3:3]) ^ (matrix1[0][2:2]&AT2in1[2:2]) ^ (matrix1[0][1:1]&AT2in1[1:1]) ^ (matrix1[0][0:0]&AT2in1[0:0]); 
assign AT2out1[6:6] = (matrix1[1][7:7]&AT2in1[7:7]) ^ (matrix1[1][6:6]&AT2in1[6:6]) ^ (matrix1[1][5:5]&AT2in1[5:5]) ^ (matrix1[1][4:4]&AT2in1[4:4]) ^ (matrix1[1][3:3]&AT2in1[3:3]) ^ (matrix1[1][2:2]&AT2in1[2:2]) ^ (matrix1[1][1:1]&AT2in1[1:1]) ^ (matrix1[1][0:0]&AT2in1[0:0]); 
assign AT2out1[5:5] = (matrix1[2][7:7]&AT2in1[7:7]) ^ (matrix1[2][6:6]&AT2in1[6:6]) ^ (matrix1[2][5:5]&AT2in1[5:5]) ^ (matrix1[2][4:4]&AT2in1[4:4]) ^ (matrix1[2][3:3]&AT2in1[3:3]) ^ (matrix1[2][2:2]&AT2in1[2:2]) ^ (matrix1[2][1:1]&AT2in1[1:1]) ^ (matrix1[2][0:0]&AT2in1[0:0]); 
assign AT2out1[4:4] = (matrix1[3][7:7]&AT2in1[7:7]) ^ (matrix1[3][6:6]&AT2in1[6:6]) ^ (matrix1[3][5:5]&AT2in1[5:5]) ^ (matrix1[3][4:4]&AT2in1[4:4]) ^ (matrix1[3][3:3]&AT2in1[3:3]) ^ (matrix1[3][2:2]&AT2in1[2:2]) ^ (matrix1[3][1:1]&AT2in1[1:1]) ^ (matrix1[3][0:0]&AT2in1[0:0]); 
assign AT2out1[3:3] = (matrix1[4][7:7]&AT2in1[7:7]) ^ (matrix1[4][6:6]&AT2in1[6:6]) ^ (matrix1[4][5:5]&AT2in1[5:5]) ^ (matrix1[4][4:4]&AT2in1[4:4]) ^ (matrix1[4][3:3]&AT2in1[3:3]) ^ (matrix1[4][2:2]&AT2in1[2:2]) ^ (matrix1[4][1:1]&AT2in1[1:1]) ^ (matrix1[4][0:0]&AT2in1[0:0]); 
assign AT2out1[2:2] = (matrix1[5][7:7]&AT2in1[7:7]) ^ (matrix1[5][6:6]&AT2in1[6:6]) ^ (matrix1[5][5:5]&AT2in1[5:5]) ^ (matrix1[5][4:4]&AT2in1[4:4]) ^ (matrix1[5][3:3]&AT2in1[3:3]) ^ (matrix1[5][2:2]&AT2in1[2:2]) ^ (matrix1[5][1:1]&AT2in1[1:1]) ^ (matrix1[5][0:0]&AT2in1[0:0]); 
assign AT2out1[1:1] = (matrix1[6][7:7]&AT2in1[7:7]) ^ (matrix1[6][6:6]&AT2in1[6:6]) ^ (matrix1[6][5:5]&AT2in1[5:5]) ^ (matrix1[6][4:4]&AT2in1[4:4]) ^ (matrix1[6][3:3]&AT2in1[3:3]) ^ (matrix1[6][2:2]&AT2in1[2:2]) ^ (matrix1[6][1:1]&AT2in1[1:1]) ^ (matrix1[6][0:0]&AT2in1[0:0]); 
assign AT2out1[0:0] = (matrix1[7][7:7]&AT2in1[7:7]) ^ (matrix1[7][6:6]&AT2in1[6:6]) ^ (matrix1[7][5:5]&AT2in1[5:5]) ^ (matrix1[7][4:4]&AT2in1[4:4]) ^ (matrix1[7][3:3]&AT2in1[3:3]) ^ (matrix1[7][2:2]&AT2in1[2:2]) ^ (matrix1[7][1:1]&AT2in1[1:1]) ^ (matrix1[7][0:0]&AT2in1[0:0]); 

assign sbout0 = AT2out0;
assign sbout1 = AT2out1;



endmodule

