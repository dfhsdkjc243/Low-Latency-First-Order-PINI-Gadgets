module Stage23_smt_trivialopt_l4_PINI(
input clk,
input [11:0] a0b0c0d0e0f0g0h0i0j0k0l0,
input [11:0] a1b1c1d1e1f1g1h1i1j1k1l1,
input [21:0] ran,
output [7:0] x0y0z0t0m0n0p0q0,
output [7:0] x1y1z1t1m1n1p1q1
);


wire a0_i,b0_i,c0_i,d0_i,e0_i,f0_i,g0_i,h0_i;
wire a1_i,b1_i,c1_i,d1_i,e1_i,f1_i,g1_i,h1_i;
wire a0,b0,c0,d0,e0,f0,g0,h0;
wire a1,b1,c1,d1,e1,f1,g1,h1;
wire x0,y0,z0,t0,m0,n0,p0,q0;
wire x1,y1,z1,t1,m1,n1,p1,q1;
wire i0,j0,k0,l0;
wire i1,j1,k1,l1;
wire r0m, r1m, r2m, r3m, r4m, r5m, r6m, r7m, r8m, r9m, r10m, r11m, r12m, r13m, r14m, r15m, r16m, r17m, r18m, r19m, r20m, r21m;

//pow4
assign {j0_i,i0_i,l0_i,k0_i,h0_i,g0_i,f0_i,e0_i,d0_i,c0_i,b0_i,a0_i} = a0b0c0d0e0f0g0h0i0j0k0l0;
assign {j1_i,i1_i,l1_i,k1_i,h1_i,g1_i,f1_i,e1_i,d1_i,c1_i,b1_i,a1_i} = a1b1c1d1e1f1g1h1i1j1k1l1;


assign {h0,g0,f0,e0,d0,c0,b0,a0} = {h0_i,g0_i,f0_i,e0_i,d0_i,c0_i,b0_i,a0_i};
assign {h1,g1,f1,e1,d1,c1,b1,a1} = {h1_i,g1_i,f1_i,e1_i,d1_i,c1_i,b1_i,a1_i};

assign	  i0 = (i0_i ^ j0_i);
assign    j0 = (j0_i ^ k0_i);
assign    k0 = (k0_i)       ;
assign    l0 = (l0_i)       ;

assign	  i1 = (i1_i ^ j1_i);
assign    j1 = (j1_i ^ k1_i);
assign    k1 = (k1_i)       ;
assign    l1 = (l1_i)       ;



assign {r0m, r1m, r2m, r3m, r4m, r5m, r6m, r7m, r8m, r9m, r10m, r11m, r12m, r13m, r14m, r15m, r16m, r17m, r18m, r19m, r20m, r21m} = ran;

reg reg_0_0, reg_0_1, reg_0_2, reg_0_3, reg_0_4, reg_0_5, reg_0_6, reg_0_7, reg_0_8, reg_0_9, reg_0_10, reg_0_11, reg_0_12, reg_0_13, reg_0_14, reg_0_15, reg_0_16, reg_0_17, reg_0_18, reg_0_19, reg_0_20, reg_0_21, reg_0_22, reg_0_23, reg_0_24, reg_0_25, reg_0_26, reg_0_27, reg_0_28, reg_0_29, reg_0_30, reg_0_31, reg_0_32, reg_0_33;
reg reg_1_0, reg_1_1, reg_1_2, reg_1_3, reg_1_4, reg_1_5, reg_1_6, reg_1_7, reg_1_8, reg_1_9, reg_1_10, reg_1_11, reg_1_12, reg_1_13, reg_1_14, reg_1_15, reg_1_16, reg_1_17, reg_1_18, reg_1_19, reg_1_20, reg_1_21, reg_1_22, reg_1_23, reg_1_24, reg_1_25, reg_1_26, reg_1_27, reg_1_28, reg_1_29, reg_1_30, reg_1_31, reg_1_32, reg_1_33;


wire cdx_0m = (i1 ^ r0m);
wire cdx_1m = (j1 ^ r1m);
wire cdx_2m = (k1 ^ r2m);
wire cdx_3m = (l1 ^ r3m);
wire cdx_4m = i1&j1 ^ r4m;
wire cdx_5m = i1&k1 ^ r5m;
wire cdx_6m = i1&l1 ^ r6m;
wire cdx_7m = j1&k1 ^ r7m;
wire cdx_8m = j1&l1 ^ r8m;
wire cdx_9m = k1&l1 ^ r9m;
wire cdx_10m = i1&j1&k1 ^ r10m;
wire cdx_11m = i1&j1&l1 ^ r11m;
wire cdx_12m = i1&k1&l1 ^ r12m;
wire cdx_13m = j1&k1&l1 ^ r13m;
wire cdx_14m = i0 ^ r0m;
wire cdx_15m = (cdx_14m);
wire cdx_16m = e0&cdx_15m;
wire cdx_17m = (reg_0_12);
wire cdx_18m = (cdx_17m);
wire cdx_19m = reg_0_4&cdx_18m;
wire cdx_20m = j0 ^ r1m;
wire cdx_21m = (cdx_20m);
wire cdx_22m = e0&cdx_21m;
wire cdx_23m = (reg_0_13);
wire cdx_24m = (cdx_23m);
wire cdx_25m = reg_0_4&cdx_24m;
wire cdx_26m = l0 ^ r3m;
wire cdx_27m = (cdx_26m);
wire cdx_28m = e0&cdx_27m;
wire cdx_29m = (reg_0_15);
wire cdx_30m = (cdx_29m);
wire cdx_31m = reg_0_4&cdx_30m;
wire cdx_32m = f0&cdx_15m;
wire cdx_33m = reg_0_5&cdx_18m;
wire cdx_34m = g0&cdx_15m;
wire cdx_35m = reg_0_6&cdx_18m;
wire cdx_36m = g0&cdx_21m;
wire cdx_37m = reg_0_6&cdx_24m;
wire cdx_38m = k0 ^ r2m;
wire cdx_39m = (cdx_38m);
wire cdx_40m = g0&cdx_39m;
wire cdx_41m = (reg_0_14);
wire cdx_42m = (cdx_41m);
wire cdx_43m = reg_0_6&cdx_42m;
wire cdx_44m = h0&cdx_15m;
wire cdx_45m = reg_0_7&cdx_18m;
wire cdx_46m = h0&cdx_39m;
wire cdx_47m = reg_0_7&cdx_42m;
wire cdx_48m = h0&cdx_27m;
wire cdx_49m = reg_0_7&cdx_30m;
wire cdx_50m = j0&k0 ^ r7m;
wire cdx_51m = k0;
wire cdx_52m = j0;
wire cdx_53m = cdx_51m&r11m;
wire cdx_54m = cdx_52m&r12m;
wire cdx_55m = (cdx_50m ^ cdx_51m&r1m ^ cdx_52m&r2m);
wire cdx_56m = e0&cdx_55m;
wire cdx_57m = (reg_0_19);
wire cdx_58m = reg_0_10&cdx_23m;
wire cdx_59m = reg_0_9&cdx_41m;
wire cdx_60m = (cdx_58m ^ cdx_59m ^ cdx_57m);
wire cdx_61m = reg_0_4&cdx_60m;
wire cdx_62m = i0&l0 ^ r6m;
wire cdx_63m = l0;
wire cdx_64m = i0;
wire cdx_65m = cdx_63m&r10m;
wire cdx_66m = cdx_64m&r13m;
wire cdx_67m = (cdx_62m ^ cdx_63m&r0m ^ cdx_64m&r3m);
wire cdx_68m = f0&cdx_67m;
wire cdx_69m = (reg_0_18);
wire cdx_70m = reg_0_11&cdx_17m;
wire cdx_71m = reg_0_8&cdx_29m;
wire cdx_72m = (cdx_70m ^ cdx_71m ^ cdx_69m);
wire cdx_73m = reg_0_5&cdx_72m;
wire cdx_74m = f0&cdx_55m;
wire cdx_75m = reg_0_5&cdx_60m;
wire cdx_76m = cdx_52m&cdx_63m ^ r8m;
wire cdx_77m = cdx_63m&r11m;
wire cdx_78m = cdx_52m&r13m;
wire cdx_79m = (cdx_76m ^ cdx_63m&r1m ^ cdx_52m&r3m);
wire cdx_80m = f0&cdx_79m;
wire cdx_81m = (reg_0_20);
wire cdx_82m = reg_0_11&cdx_23m;
wire cdx_83m = reg_0_9&cdx_29m;
wire cdx_84m = (cdx_82m ^ cdx_83m ^ cdx_81m);
wire cdx_85m = reg_0_5&cdx_84m;
wire cdx_86m = g0&cdx_67m;
wire cdx_87m = reg_0_6&cdx_72m;
wire cdx_88m = g0&cdx_55m;
wire cdx_89m = reg_0_6&cdx_60m;
wire cdx_90m = cdx_51m&cdx_63m ^ r9m;
wire cdx_91m = cdx_63m&r12m;
wire cdx_92m = cdx_51m&r13m;
wire cdx_93m = (cdx_90m ^ cdx_63m&r2m ^ cdx_51m&r3m);
wire cdx_94m = g0&cdx_93m;
wire cdx_95m = (reg_0_21);
wire cdx_96m = reg_0_11&cdx_41m;
wire cdx_97m = reg_0_10&cdx_29m;
wire cdx_98m = (cdx_96m ^ cdx_97m ^ cdx_95m);
wire cdx_99m = reg_0_6&cdx_98m;
wire cdx_100m = cdx_64m&cdx_51m ^ r5m;
wire cdx_101m = cdx_51m&r10m;
wire cdx_102m = cdx_64m&r12m;
wire cdx_103m = (cdx_100m ^ cdx_51m&r0m ^ cdx_64m&r2m);
wire cdx_104m = h0&cdx_103m;
wire cdx_105m = (reg_0_17);
wire cdx_106m = reg_0_10&cdx_17m;
wire cdx_107m = reg_0_8&cdx_41m;
wire cdx_108m = (cdx_106m ^ cdx_107m ^ cdx_105m);
wire cdx_109m = reg_0_7&cdx_108m;
wire cdx_110m = h0&cdx_67m;
wire cdx_111m = reg_0_7&cdx_72m;
wire cdx_112m = h0&cdx_79m;
wire cdx_113m = reg_0_7&cdx_84m;
wire cdx_114m = cdx_64m&cdx_52m&cdx_63m ^ r11m;
wire cdx_115m = cdx_52m&cdx_63m;
wire cdx_116m = cdx_64m&cdx_63m;
wire cdx_117m = cdx_64m&cdx_52m;
wire cdx_118m = cdx_52m&cdx_65m;
wire cdx_119m = cdx_64m&cdx_77m;
wire cdx_120m = cdx_64m&cdx_78m;
wire cdx_121m = cdx_63m&r0m;
wire cdx_122m = cdx_52m&r2m;
wire cdx_123m = cdx_64m&r4m;
wire cdx_124m = (cdx_114m ^ cdx_115m&r0m ^ cdx_116m&r1m ^ cdx_117m&r3m ^ cdx_63m&r4m ^ cdx_52m&r6m ^ cdx_64m&r8m);
wire cdx_125m = e0&cdx_124m;
wire cdx_126m = (reg_0_16);
wire cdx_127m = (reg_0_23);
wire cdx_128m = reg_0_9&cdx_70m;
wire cdx_129m = reg_0_8&cdx_82m;
wire cdx_130m = reg_0_8&cdx_83m;
wire cdx_131m = reg_0_11&cdx_126m;
wire cdx_132m = reg_0_9&cdx_69m;
wire cdx_133m = reg_0_8&cdx_81m;
wire cdx_134m = (cdx_128m ^ cdx_129m ^ cdx_130m ^ cdx_131m ^ cdx_132m ^ cdx_133m ^ cdx_127m);
wire cdx_135m = reg_0_4&cdx_134m;
wire cdx_136m = cdx_117m&cdx_51m ^ r10m;
wire cdx_137m = cdx_52m&cdx_51m;
wire cdx_138m = cdx_64m&cdx_51m;
wire cdx_139m = cdx_52m&cdx_101m;
wire cdx_140m = cdx_64m&cdx_53m;
wire cdx_141m = cdx_64m&cdx_54m;
wire cdx_142m = cdx_51m&r0m;
wire cdx_143m = cdx_52m&r1m;
wire cdx_144m = cdx_64m&r3m;
wire cdx_145m = (cdx_136m ^ cdx_137m&r0m ^ cdx_138m&r1m ^ cdx_117m&r2m ^ cdx_51m&r4m ^ cdx_52m&r5m ^ cdx_64m&r7m);
wire cdx_146m = f0&cdx_145m;
wire cdx_147m = (reg_0_22);
wire cdx_148m = reg_0_9&cdx_106m;
wire cdx_149m = reg_0_8&cdx_58m;
wire cdx_150m = reg_0_8&cdx_59m;
wire cdx_151m = reg_0_10&cdx_126m;
wire cdx_152m = reg_0_9&cdx_105m;
wire cdx_153m = reg_0_8&cdx_57m;
wire cdx_154m = (cdx_148m ^ cdx_149m ^ cdx_150m ^ cdx_151m ^ cdx_152m ^ cdx_153m ^ cdx_147m);
wire cdx_155m = reg_0_5&cdx_154m;
wire cdx_156m = cdx_137m&cdx_63m ^ r13m;
wire cdx_157m = cdx_51m&cdx_63m;
wire cdx_158m = cdx_51m&cdx_77m;
wire cdx_159m = cdx_52m&cdx_91m;
wire cdx_160m = cdx_52m&cdx_92m;
wire cdx_161m = cdx_63m&r3m;
wire cdx_162m = cdx_51m&r4m;
wire cdx_163m = cdx_52m&r5m;
wire cdx_164m = (cdx_156m ^ cdx_157m&r1m ^ cdx_115m&r2m ^ cdx_137m&r3m ^ cdx_63m&r7m ^ cdx_51m&r8m ^ cdx_52m&r9m);
wire cdx_165m = f0&cdx_164m;
wire cdx_166m = (reg_0_25);
wire cdx_167m = reg_0_10&cdx_82m;
wire cdx_168m = reg_0_9&cdx_96m;
wire cdx_169m = reg_0_9&cdx_97m;
wire cdx_170m = reg_0_11&cdx_57m;
wire cdx_171m = reg_0_10&cdx_81m;
wire cdx_172m = reg_0_9&cdx_95m;
wire cdx_173m = (cdx_167m ^ cdx_168m ^ cdx_169m ^ cdx_170m ^ cdx_171m ^ cdx_172m ^ cdx_166m);
wire cdx_174m = reg_0_5&cdx_173m;
wire cdx_175m = g0&cdx_124m;
wire cdx_176m = reg_0_6&cdx_134m;
wire cdx_177m = cdx_138m&cdx_63m ^ r12m;
wire cdx_178m = cdx_51m&cdx_65m;
wire cdx_179m = cdx_64m&cdx_91m;
wire cdx_180m = cdx_64m&cdx_92m;
wire cdx_181m = cdx_63m&r1m;
wire cdx_182m = cdx_51m&r2m;
wire cdx_183m = cdx_64m&r5m;
wire cdx_184m = (cdx_177m ^ cdx_51m&cdx_121m ^ cdx_116m&r2m ^ cdx_138m&r3m ^ cdx_63m&r5m ^ cdx_51m&r6m ^ cdx_64m&r9m);
wire cdx_185m = g0&cdx_184m;
wire cdx_186m = (reg_0_24);
wire cdx_187m = reg_0_10&cdx_70m;
wire cdx_188m = reg_0_8&cdx_96m;
wire cdx_189m = reg_0_8&cdx_97m;
wire cdx_190m = reg_0_11&cdx_105m;
wire cdx_191m = reg_0_10&cdx_69m;
wire cdx_192m = reg_0_8&cdx_95m;
wire cdx_193m = (cdx_187m ^ cdx_188m ^ cdx_189m ^ cdx_190m ^ cdx_191m ^ cdx_192m ^ cdx_186m);
wire cdx_194m = reg_0_6&cdx_193m;
wire cdx_195m = g0&cdx_164m;
wire cdx_196m = reg_0_6&cdx_173m;
wire cdx_197m = h0&cdx_145m;
wire cdx_198m = reg_0_7&cdx_154m;
wire cdx_199m = h0&cdx_184m;
wire cdx_200m = reg_0_7&cdx_193m;
wire cdx_201m = h0&cdx_164m;
wire cdx_202m = reg_0_7&cdx_173m;
wire cdx_203m = f0&cdx_21m;
wire cdx_204m = reg_0_5&cdx_24m;
wire cdx_205m = f0&cdx_27m;
wire cdx_206m = reg_0_5&cdx_30m;
wire cdx_207m = g0&cdx_27m;
wire cdx_208m = reg_0_6&cdx_30m;
wire cdx_209m = h0&cdx_21m;
wire cdx_210m = reg_0_7&cdx_24m;
wire cdx_211m = e0&cdx_67m;
wire cdx_212m = reg_0_4&cdx_72m;
wire cdx_213m = e0&cdx_79m;
wire cdx_214m = reg_0_4&cdx_84m;
wire cdx_215m = g0&cdx_103m;
wire cdx_216m = reg_0_6&cdx_108m;
wire cdx_217m = g0&cdx_79m;
wire cdx_218m = reg_0_6&cdx_84m;
wire cdx_219m = h0&cdx_55m;
wire cdx_220m = reg_0_7&cdx_60m;
wire cdx_221m = h0&cdx_93m;
wire cdx_222m = reg_0_7&cdx_98m;
wire cdx_223m = e0&cdx_145m;
wire cdx_224m = reg_0_4&cdx_154m;
wire cdx_225m = e0&cdx_164m;
wire cdx_226m = reg_0_4&cdx_173m;
wire cdx_227m = f0&cdx_124m;
wire cdx_228m = reg_0_5&cdx_134m;
wire cdx_229m = g0&cdx_145m;
wire cdx_230m = reg_0_6&cdx_154m;
wire cdx_231m = h0&cdx_124m;
wire cdx_232m = reg_0_7&cdx_134m;
wire cdx_233m = e0&cdx_39m;
wire cdx_234m = reg_0_4&cdx_42m;
wire cdx_235m = f0&cdx_39m;
wire cdx_236m = reg_0_5&cdx_42m;
wire cdx_237m = e0&cdx_93m;
wire cdx_238m = reg_0_4&cdx_98m;
wire cdx_239m = f0&cdx_103m;
wire cdx_240m = reg_0_5&cdx_108m;
wire cdx_241m = e0&cdx_184m;
wire cdx_242m = reg_0_4&cdx_193m;
wire cdx_243m = f0&cdx_184m;
wire cdx_244m = reg_0_5&cdx_193m;
wire cdx_245m = e0&cdx_103m;
wire cdx_246m = reg_0_4&cdx_108m;
wire cdx_247m = f0&cdx_93m;
wire cdx_248m = reg_0_5&cdx_98m;
wire cdx_249m = a0&cdx_15m;
wire cdx_250m = reg_0_0&cdx_18m;
wire cdx_251m = a0&cdx_21m;
wire cdx_252m = reg_0_0&cdx_24m;
wire cdx_253m = a0&cdx_27m;
wire cdx_254m = reg_0_0&cdx_30m;
wire cdx_255m = b0&cdx_15m;
wire cdx_256m = reg_0_1&cdx_18m;
wire cdx_257m = c0&cdx_15m;
wire cdx_258m = reg_0_2&cdx_18m;
wire cdx_259m = c0&cdx_21m;
wire cdx_260m = reg_0_2&cdx_24m;
wire cdx_261m = c0&cdx_39m;
wire cdx_262m = reg_0_2&cdx_42m;
wire cdx_263m = d0&cdx_15m;
wire cdx_264m = reg_0_3&cdx_18m;
wire cdx_265m = d0&cdx_39m;
wire cdx_266m = reg_0_3&cdx_42m;
wire cdx_267m = d0&cdx_27m;
wire cdx_268m = reg_0_3&cdx_30m;
wire cdx_269m = a0&cdx_55m;
wire cdx_270m = reg_0_0&cdx_60m;
wire cdx_271m = b0&cdx_67m;
wire cdx_272m = reg_0_1&cdx_72m;
wire cdx_273m = b0&cdx_55m;
wire cdx_274m = reg_0_1&cdx_60m;
wire cdx_275m = b0&cdx_79m;
wire cdx_276m = reg_0_1&cdx_84m;
wire cdx_277m = c0&cdx_67m;
wire cdx_278m = reg_0_2&cdx_72m;
wire cdx_279m = c0&cdx_55m;
wire cdx_280m = reg_0_2&cdx_60m;
wire cdx_281m = c0&cdx_93m;
wire cdx_282m = reg_0_2&cdx_98m;
wire cdx_283m = d0&cdx_103m;
wire cdx_284m = reg_0_3&cdx_108m;
wire cdx_285m = d0&cdx_67m;
wire cdx_286m = reg_0_3&cdx_72m;
wire cdx_287m = d0&cdx_79m;
wire cdx_288m = reg_0_3&cdx_84m;
wire cdx_289m = a0&cdx_124m;
wire cdx_290m = reg_0_0&cdx_134m;
wire cdx_291m = b0&cdx_145m;
wire cdx_292m = reg_0_1&cdx_154m;
wire cdx_293m = b0&cdx_164m;
wire cdx_294m = reg_0_1&cdx_173m;
wire cdx_295m = c0&cdx_124m;
wire cdx_296m = reg_0_2&cdx_134m;
wire cdx_297m = c0&cdx_184m;
wire cdx_298m = reg_0_2&cdx_193m;
wire cdx_299m = c0&cdx_164m;
wire cdx_300m = reg_0_2&cdx_173m;
wire cdx_301m = d0&cdx_145m;
wire cdx_302m = reg_0_3&cdx_154m;
wire cdx_303m = d0&cdx_184m;
wire cdx_304m = reg_0_3&cdx_193m;
wire cdx_305m = d0&cdx_164m;
wire cdx_306m = reg_0_3&cdx_173m;
wire cdx_307m = b0&cdx_21m;
wire cdx_308m = reg_0_1&cdx_24m;
wire cdx_309m = b0&cdx_27m;
wire cdx_310m = reg_0_1&cdx_30m;
wire cdx_311m = c0&cdx_27m;
wire cdx_312m = reg_0_2&cdx_30m;
wire cdx_313m = d0&cdx_21m;
wire cdx_314m = reg_0_3&cdx_24m;
wire cdx_315m = a0&cdx_67m;
wire cdx_316m = reg_0_0&cdx_72m;
wire cdx_317m = a0&cdx_79m;
wire cdx_318m = reg_0_0&cdx_84m;
wire cdx_319m = c0&cdx_103m;
wire cdx_320m = reg_0_2&cdx_108m;
wire cdx_321m = c0&cdx_79m;
wire cdx_322m = reg_0_2&cdx_84m;
wire cdx_323m = d0&cdx_55m;
wire cdx_324m = reg_0_3&cdx_60m;
wire cdx_325m = d0&cdx_93m;
wire cdx_326m = reg_0_3&cdx_98m;
wire cdx_327m = a0&cdx_145m;
wire cdx_328m = reg_0_0&cdx_154m;
wire cdx_329m = a0&cdx_164m;
wire cdx_330m = reg_0_0&cdx_173m;
wire cdx_331m = b0&cdx_124m;
wire cdx_332m = reg_0_1&cdx_134m;
wire cdx_333m = c0&cdx_145m;
wire cdx_334m = reg_0_2&cdx_154m;
wire cdx_335m = d0&cdx_124m;
wire cdx_336m = reg_0_3&cdx_134m;
wire cdx_337m = a0&cdx_39m;
wire cdx_338m = reg_0_0&cdx_42m;
wire cdx_339m = b0&cdx_39m;
wire cdx_340m = reg_0_1&cdx_42m;
wire cdx_341m = a0&cdx_93m;
wire cdx_342m = reg_0_0&cdx_98m;
wire cdx_343m = b0&cdx_103m;
wire cdx_344m = reg_0_1&cdx_108m;
wire cdx_345m = a0&cdx_184m;
wire cdx_346m = reg_0_0&cdx_193m;
wire cdx_347m = b0&cdx_184m;
wire cdx_348m = reg_0_1&cdx_193m;
wire cdx_349m = a0&cdx_103m;
wire cdx_350m = reg_0_0&cdx_108m;
wire cdx_351m = b0&cdx_93m;
wire cdx_352m = reg_0_1&cdx_98m;
wire cdx_353m = cdx_117m ^ r4m;
wire cdx_354m = i1 ^ r0m;
wire cdx_355m = e1&cdx_0m;
wire cdx_356m = (reg_1_12);
wire cdx_357m = (cdx_356m);
wire cdx_358m = reg_1_4&cdx_357m;
wire cdx_359m = j1 ^ r1m;
wire cdx_360m = e1&cdx_1m;
wire cdx_361m = (reg_1_13);
wire cdx_362m = (cdx_361m);
wire cdx_363m = reg_1_4&cdx_362m;
wire cdx_364m = l1 ^ r3m;
wire cdx_365m = e1&cdx_3m;
wire cdx_366m = (reg_1_15);
wire cdx_367m = (cdx_366m);
wire cdx_368m = reg_1_4&cdx_367m;
wire cdx_369m = f1&cdx_0m;
wire cdx_370m = reg_1_5&cdx_357m;
wire cdx_371m = g1&cdx_0m;
wire cdx_372m = reg_1_6&cdx_357m;
wire cdx_373m = g1&cdx_1m;
wire cdx_374m = reg_1_6&cdx_362m;
wire cdx_375m = k1 ^ r2m;
wire cdx_376m = g1&cdx_2m;
wire cdx_377m = (reg_1_14);
wire cdx_378m = (cdx_377m);
wire cdx_379m = reg_1_6&cdx_378m;
wire cdx_380m = h1&cdx_0m;
wire cdx_381m = reg_1_7&cdx_357m;
wire cdx_382m = h1&cdx_2m;
wire cdx_383m = reg_1_7&cdx_378m;
wire cdx_384m = h1&cdx_3m;
wire cdx_385m = reg_1_7&cdx_367m;
wire cdx_386m = k1;
wire cdx_387m = j1;
wire cdx_388m = cdx_386m&r11m;
wire cdx_389m = cdx_387m&r12m;
wire cdx_390m = (cdx_7m ^ cdx_386m&r1m ^ cdx_387m&r2m);
wire cdx_391m = e1&cdx_390m;
wire cdx_392m = (reg_1_19);
wire cdx_393m = reg_1_10&cdx_361m;
wire cdx_394m = reg_1_9&cdx_377m;
wire cdx_395m = (cdx_393m ^ cdx_394m ^ cdx_392m);
wire cdx_396m = reg_1_4&cdx_395m;
wire cdx_397m = l1;
wire cdx_398m = i1;
wire cdx_399m = cdx_397m&r10m;
wire cdx_400m = cdx_398m&r13m;
wire cdx_401m = (cdx_6m ^ cdx_397m&r0m ^ cdx_398m&r3m);
wire cdx_402m = f1&cdx_401m;
wire cdx_403m = (reg_1_18);
wire cdx_404m = reg_1_11&cdx_356m;
wire cdx_405m = reg_1_8&cdx_366m;
wire cdx_406m = (cdx_404m ^ cdx_405m ^ cdx_403m);
wire cdx_407m = reg_1_5&cdx_406m;
wire cdx_408m = f1&cdx_390m;
wire cdx_409m = reg_1_5&cdx_395m;
wire cdx_410m = cdx_397m&r11m;
wire cdx_411m = cdx_387m&r13m;
wire cdx_412m = (cdx_8m ^ cdx_397m&r1m ^ cdx_387m&r3m);
wire cdx_413m = f1&cdx_412m;
wire cdx_414m = (reg_1_20);
wire cdx_415m = reg_1_11&cdx_361m;
wire cdx_416m = reg_1_9&cdx_366m;
wire cdx_417m = (cdx_415m ^ cdx_416m ^ cdx_414m);
wire cdx_418m = reg_1_5&cdx_417m;
wire cdx_419m = g1&cdx_401m;
wire cdx_420m = reg_1_6&cdx_406m;
wire cdx_421m = g1&cdx_390m;
wire cdx_422m = reg_1_6&cdx_395m;
wire cdx_423m = cdx_397m&r12m;
wire cdx_424m = cdx_386m&r13m;
wire cdx_425m = (cdx_9m ^ cdx_397m&r2m ^ cdx_386m&r3m);
wire cdx_426m = g1&cdx_425m;
wire cdx_427m = (reg_1_21);
wire cdx_428m = reg_1_11&cdx_377m;
wire cdx_429m = reg_1_10&cdx_366m;
wire cdx_430m = (cdx_428m ^ cdx_429m ^ cdx_427m);
wire cdx_431m = reg_1_6&cdx_430m;
wire cdx_432m = cdx_386m&r10m;
wire cdx_433m = cdx_398m&r12m;
wire cdx_434m = (cdx_5m ^ cdx_386m&r0m ^ cdx_398m&r2m);
wire cdx_435m = h1&cdx_434m;
wire cdx_436m = (reg_1_17);
wire cdx_437m = reg_1_10&cdx_356m;
wire cdx_438m = reg_1_8&cdx_377m;
wire cdx_439m = (cdx_437m ^ cdx_438m ^ cdx_436m);
wire cdx_440m = reg_1_7&cdx_439m;
wire cdx_441m = h1&cdx_401m;
wire cdx_442m = reg_1_7&cdx_406m;
wire cdx_443m = h1&cdx_412m;
wire cdx_444m = reg_1_7&cdx_417m;
wire cdx_445m = cdx_387m&cdx_397m;
wire cdx_446m = cdx_398m&cdx_397m;
wire cdx_447m = cdx_398m&cdx_387m;
wire cdx_448m = cdx_387m&cdx_399m;
wire cdx_449m = cdx_398m&cdx_410m;
wire cdx_450m = cdx_398m&cdx_411m;
wire cdx_451m = cdx_397m&r0m;
wire cdx_452m = cdx_387m&r2m;
wire cdx_453m = cdx_398m&r4m;
wire cdx_454m = (cdx_11m ^ cdx_445m&r0m ^ cdx_446m&r1m ^ cdx_447m&r3m ^ cdx_397m&r4m ^ cdx_387m&r6m ^ cdx_398m&r8m);
wire cdx_455m = e1&cdx_454m;
wire cdx_456m = (reg_1_16);
wire cdx_457m = (reg_1_23);
wire cdx_458m = reg_1_9&cdx_404m;
wire cdx_459m = reg_1_8&cdx_415m;
wire cdx_460m = reg_1_8&cdx_416m;
wire cdx_461m = reg_1_11&cdx_456m;
wire cdx_462m = reg_1_9&cdx_403m;
wire cdx_463m = reg_1_8&cdx_414m;
wire cdx_464m = (cdx_458m ^ cdx_459m ^ cdx_460m ^ cdx_461m ^ cdx_462m ^ cdx_463m ^ cdx_457m);
wire cdx_465m = reg_1_4&cdx_464m;
wire cdx_466m = cdx_387m&cdx_386m;
wire cdx_467m = cdx_398m&cdx_386m;
wire cdx_468m = cdx_387m&cdx_432m;
wire cdx_469m = cdx_398m&cdx_388m;
wire cdx_470m = cdx_398m&cdx_389m;
wire cdx_471m = cdx_386m&r0m;
wire cdx_472m = cdx_387m&r1m;
wire cdx_473m = cdx_398m&r3m;
wire cdx_474m = (cdx_10m ^ cdx_466m&r0m ^ cdx_467m&r1m ^ cdx_447m&r2m ^ cdx_386m&r4m ^ cdx_387m&r5m ^ cdx_398m&r7m);
wire cdx_475m = f1&cdx_474m;
wire cdx_476m = (reg_1_22);
wire cdx_477m = reg_1_9&cdx_437m;
wire cdx_478m = reg_1_8&cdx_393m;
wire cdx_479m = reg_1_8&cdx_394m;
wire cdx_480m = reg_1_10&cdx_456m;
wire cdx_481m = reg_1_9&cdx_436m;
wire cdx_482m = reg_1_8&cdx_392m;
wire cdx_483m = (cdx_477m ^ cdx_478m ^ cdx_479m ^ cdx_480m ^ cdx_481m ^ cdx_482m ^ cdx_476m);
wire cdx_484m = reg_1_5&cdx_483m;
wire cdx_485m = cdx_386m&cdx_397m;
wire cdx_486m = cdx_386m&cdx_410m;
wire cdx_487m = cdx_387m&cdx_423m;
wire cdx_488m = cdx_387m&cdx_424m;
wire cdx_489m = cdx_397m&r3m;
wire cdx_490m = cdx_386m&r4m;
wire cdx_491m = cdx_387m&r5m;
wire cdx_492m = (cdx_13m ^ cdx_485m&r1m ^ cdx_445m&r2m ^ cdx_466m&r3m ^ cdx_397m&r7m ^ cdx_386m&r8m ^ cdx_387m&r9m);
wire cdx_493m = f1&cdx_492m;
wire cdx_494m = (reg_1_25);
wire cdx_495m = reg_1_10&cdx_415m;
wire cdx_496m = reg_1_9&cdx_428m;
wire cdx_497m = reg_1_9&cdx_429m;
wire cdx_498m = reg_1_11&cdx_392m;
wire cdx_499m = reg_1_10&cdx_414m;
wire cdx_500m = reg_1_9&cdx_427m;
wire cdx_501m = (cdx_495m ^ cdx_496m ^ cdx_497m ^ cdx_498m ^ cdx_499m ^ cdx_500m ^ cdx_494m);
wire cdx_502m = reg_1_5&cdx_501m;
wire cdx_503m = g1&cdx_454m;
wire cdx_504m = reg_1_6&cdx_464m;
wire cdx_505m = cdx_386m&cdx_399m;
wire cdx_506m = cdx_398m&cdx_423m;
wire cdx_507m = cdx_398m&cdx_424m;
wire cdx_508m = cdx_397m&r1m;
wire cdx_509m = cdx_386m&r2m;
wire cdx_510m = cdx_398m&r5m;
wire cdx_511m = (cdx_12m ^ cdx_386m&cdx_451m ^ cdx_446m&r2m ^ cdx_467m&r3m ^ cdx_397m&r5m ^ cdx_386m&r6m ^ cdx_398m&r9m);
wire cdx_512m = g1&cdx_511m;
wire cdx_513m = (reg_1_24);
wire cdx_514m = reg_1_10&cdx_404m;
wire cdx_515m = reg_1_8&cdx_428m;
wire cdx_516m = reg_1_8&cdx_429m;
wire cdx_517m = reg_1_11&cdx_436m;
wire cdx_518m = reg_1_10&cdx_403m;
wire cdx_519m = reg_1_8&cdx_427m;
wire cdx_520m = (cdx_514m ^ cdx_515m ^ cdx_516m ^ cdx_517m ^ cdx_518m ^ cdx_519m ^ cdx_513m);
wire cdx_521m = reg_1_6&cdx_520m;
wire cdx_522m = g1&cdx_492m;
wire cdx_523m = reg_1_6&cdx_501m;
wire cdx_524m = h1&cdx_474m;
wire cdx_525m = reg_1_7&cdx_483m;
wire cdx_526m = h1&cdx_511m;
wire cdx_527m = reg_1_7&cdx_520m;
wire cdx_528m = h1&cdx_492m;
wire cdx_529m = reg_1_7&cdx_501m;
wire cdx_530m = f1&cdx_1m;
wire cdx_531m = reg_1_5&cdx_362m;
wire cdx_532m = f1&cdx_3m;
wire cdx_533m = reg_1_5&cdx_367m;
wire cdx_534m = g1&cdx_3m;
wire cdx_535m = reg_1_6&cdx_367m;
wire cdx_536m = h1&cdx_1m;
wire cdx_537m = reg_1_7&cdx_362m;
wire cdx_538m = e1&cdx_401m;
wire cdx_539m = reg_1_4&cdx_406m;
wire cdx_540m = e1&cdx_412m;
wire cdx_541m = reg_1_4&cdx_417m;
wire cdx_542m = g1&cdx_434m;
wire cdx_543m = reg_1_6&cdx_439m;
wire cdx_544m = g1&cdx_412m;
wire cdx_545m = reg_1_6&cdx_417m;
wire cdx_546m = h1&cdx_390m;
wire cdx_547m = reg_1_7&cdx_395m;
wire cdx_548m = h1&cdx_425m;
wire cdx_549m = reg_1_7&cdx_430m;
wire cdx_550m = e1&cdx_474m;
wire cdx_551m = reg_1_4&cdx_483m;
wire cdx_552m = e1&cdx_492m;
wire cdx_553m = reg_1_4&cdx_501m;
wire cdx_554m = f1&cdx_454m;
wire cdx_555m = reg_1_5&cdx_464m;
wire cdx_556m = g1&cdx_474m;
wire cdx_557m = reg_1_6&cdx_483m;
wire cdx_558m = h1&cdx_454m;
wire cdx_559m = reg_1_7&cdx_464m;
wire cdx_560m = e1&cdx_2m;
wire cdx_561m = reg_1_4&cdx_378m;
wire cdx_562m = f1&cdx_2m;
wire cdx_563m = reg_1_5&cdx_378m;
wire cdx_564m = e1&cdx_425m;
wire cdx_565m = reg_1_4&cdx_430m;
wire cdx_566m = f1&cdx_434m;
wire cdx_567m = reg_1_5&cdx_439m;
wire cdx_568m = e1&cdx_511m;
wire cdx_569m = reg_1_4&cdx_520m;
wire cdx_570m = f1&cdx_511m;
wire cdx_571m = reg_1_5&cdx_520m;
wire cdx_572m = e1&cdx_434m;
wire cdx_573m = reg_1_4&cdx_439m;
wire cdx_574m = f1&cdx_425m;
wire cdx_575m = reg_1_5&cdx_430m;
wire cdx_576m = a1&cdx_0m;
wire cdx_577m = reg_1_0&cdx_357m;
wire cdx_578m = a1&cdx_1m;
wire cdx_579m = reg_1_0&cdx_362m;
wire cdx_580m = a1&cdx_3m;
wire cdx_581m = reg_1_0&cdx_367m;
wire cdx_582m = b1&cdx_0m;
wire cdx_583m = reg_1_1&cdx_357m;
wire cdx_584m = c1&cdx_0m;
wire cdx_585m = reg_1_2&cdx_357m;
wire cdx_586m = c1&cdx_1m;
wire cdx_587m = reg_1_2&cdx_362m;
wire cdx_588m = c1&cdx_2m;
wire cdx_589m = reg_1_2&cdx_378m;
wire cdx_590m = d1&cdx_0m;
wire cdx_591m = reg_1_3&cdx_357m;
wire cdx_592m = d1&cdx_2m;
wire cdx_593m = reg_1_3&cdx_378m;
wire cdx_594m = d1&cdx_3m;
wire cdx_595m = reg_1_3&cdx_367m;
wire cdx_596m = a1&cdx_390m;
wire cdx_597m = reg_1_0&cdx_395m;
wire cdx_598m = b1&cdx_401m;
wire cdx_599m = reg_1_1&cdx_406m;
wire cdx_600m = b1&cdx_390m;
wire cdx_601m = reg_1_1&cdx_395m;
wire cdx_602m = b1&cdx_412m;
wire cdx_603m = reg_1_1&cdx_417m;
wire cdx_604m = c1&cdx_401m;
wire cdx_605m = reg_1_2&cdx_406m;
wire cdx_606m = c1&cdx_390m;
wire cdx_607m = reg_1_2&cdx_395m;
wire cdx_608m = c1&cdx_425m;
wire cdx_609m = reg_1_2&cdx_430m;
wire cdx_610m = d1&cdx_434m;
wire cdx_611m = reg_1_3&cdx_439m;
wire cdx_612m = d1&cdx_401m;
wire cdx_613m = reg_1_3&cdx_406m;
wire cdx_614m = d1&cdx_412m;
wire cdx_615m = reg_1_3&cdx_417m;
wire cdx_616m = a1&cdx_454m;
wire cdx_617m = reg_1_0&cdx_464m;
wire cdx_618m = b1&cdx_474m;
wire cdx_619m = reg_1_1&cdx_483m;
wire cdx_620m = b1&cdx_492m;
wire cdx_621m = reg_1_1&cdx_501m;
wire cdx_622m = c1&cdx_454m;
wire cdx_623m = reg_1_2&cdx_464m;
wire cdx_624m = c1&cdx_511m;
wire cdx_625m = reg_1_2&cdx_520m;
wire cdx_626m = c1&cdx_492m;
wire cdx_627m = reg_1_2&cdx_501m;
wire cdx_628m = d1&cdx_474m;
wire cdx_629m = reg_1_3&cdx_483m;
wire cdx_630m = d1&cdx_511m;
wire cdx_631m = reg_1_3&cdx_520m;
wire cdx_632m = d1&cdx_492m;
wire cdx_633m = reg_1_3&cdx_501m;
wire cdx_634m = b1&cdx_1m;
wire cdx_635m = reg_1_1&cdx_362m;
wire cdx_636m = b1&cdx_3m;
wire cdx_637m = reg_1_1&cdx_367m;
wire cdx_638m = c1&cdx_3m;
wire cdx_639m = reg_1_2&cdx_367m;
wire cdx_640m = d1&cdx_1m;
wire cdx_641m = reg_1_3&cdx_362m;
wire cdx_642m = a1&cdx_401m;
wire cdx_643m = reg_1_0&cdx_406m;
wire cdx_644m = a1&cdx_412m;
wire cdx_645m = reg_1_0&cdx_417m;
wire cdx_646m = c1&cdx_434m;
wire cdx_647m = reg_1_2&cdx_439m;
wire cdx_648m = c1&cdx_412m;
wire cdx_649m = reg_1_2&cdx_417m;
wire cdx_650m = d1&cdx_390m;
wire cdx_651m = reg_1_3&cdx_395m;
wire cdx_652m = d1&cdx_425m;
wire cdx_653m = reg_1_3&cdx_430m;
wire cdx_654m = a1&cdx_474m;
wire cdx_655m = reg_1_0&cdx_483m;
wire cdx_656m = a1&cdx_492m;
wire cdx_657m = reg_1_0&cdx_501m;
wire cdx_658m = b1&cdx_454m;
wire cdx_659m = reg_1_1&cdx_464m;
wire cdx_660m = c1&cdx_474m;
wire cdx_661m = reg_1_2&cdx_483m;
wire cdx_662m = d1&cdx_454m;
wire cdx_663m = reg_1_3&cdx_464m;
wire cdx_664m = a1&cdx_2m;
wire cdx_665m = reg_1_0&cdx_378m;
wire cdx_666m = b1&cdx_2m;
wire cdx_667m = reg_1_1&cdx_378m;
wire cdx_668m = a1&cdx_425m;
wire cdx_669m = reg_1_0&cdx_430m;
wire cdx_670m = b1&cdx_434m;
wire cdx_671m = reg_1_1&cdx_439m;
wire cdx_672m = a1&cdx_511m;
wire cdx_673m = reg_1_0&cdx_520m;
wire cdx_674m = b1&cdx_511m;
wire cdx_675m = reg_1_1&cdx_520m;
wire cdx_676m = a1&cdx_434m;
wire cdx_677m = reg_1_0&cdx_439m;
wire cdx_678m = b1&cdx_425m;
wire cdx_679m = reg_1_1&cdx_430m;



always @(posedge clk) begin
	reg_0_0 <= a0;
	reg_0_1 <= b0;
	reg_0_2 <= c0;
	reg_0_3 <= d0;
	reg_0_4 <= e0;
	reg_0_5 <= f0;
	reg_0_6 <= g0;
	reg_0_7 <= h0;
	reg_0_8 <= cdx_64m;
	reg_0_9 <= cdx_52m;
	reg_0_10 <= cdx_51m;
	reg_0_11 <= cdx_63m;
	reg_0_12 <= cdx_0m;
	reg_0_13 <= cdx_1m;
	reg_0_14 <= cdx_2m;
	reg_0_15 <= cdx_3m;
	reg_0_16 <= cdx_4m;
	reg_0_17 <= cdx_5m;
	reg_0_18 <= cdx_6m;
	reg_0_19 <= cdx_7m;
	reg_0_20 <= cdx_8m;
	reg_0_21 <= cdx_9m;
	reg_0_22 <= cdx_10m;
	reg_0_23 <= cdx_11m;
	reg_0_24 <= cdx_12m;
	reg_0_25 <= cdx_13m;
	reg_0_26 <= cdx_16m ^ cdx_22m ^ cdx_28m ^ cdx_32m ^ cdx_34m ^ cdx_36m ^ cdx_40m ^ cdx_44m ^ cdx_46m ^ cdx_48m ^ cdx_56m ^ cdx_68m ^ cdx_74m ^ cdx_80m ^ cdx_86m ^ cdx_88m ^ cdx_94m ^ cdx_104m ^ cdx_110m ^ cdx_112m ^ cdx_125m ^ cdx_146m ^ cdx_165m ^ cdx_175m ^ cdx_185m ^ cdx_195m ^ cdx_197m ^ cdx_199m ^ cdx_201m ^ r14m;
	reg_0_27 <= cdx_16m ^ cdx_203m ^ cdx_205m ^ cdx_34m ^ cdx_40m ^ cdx_207m ^ cdx_209m ^ cdx_48m ^ cdx_211m ^ cdx_56m ^ cdx_213m ^ cdx_68m ^ cdx_80m ^ cdx_215m ^ cdx_86m ^ cdx_217m ^ cdx_104m ^ cdx_219m ^ cdx_112m ^ cdx_221m ^ cdx_223m ^ cdx_225m ^ cdx_146m ^ cdx_227m ^ cdx_165m ^ cdx_229m ^ cdx_185m ^ cdx_195m ^ cdx_197m ^ cdx_231m ^ r15m;
	reg_0_28 <= cdx_16m ^ cdx_22m ^ cdx_233m ^ cdx_32m ^ cdx_235m ^ cdx_205m ^ cdx_36m ^ cdx_40m ^ cdx_44m ^ cdx_209m ^ cdx_48m ^ cdx_211m ^ cdx_56m ^ cdx_237m ^ cdx_239m ^ cdx_68m ^ cdx_80m ^ cdx_215m ^ cdx_86m ^ cdx_88m ^ cdx_217m ^ cdx_104m ^ cdx_110m ^ cdx_221m ^ cdx_125m ^ cdx_241m ^ cdx_225m ^ cdx_146m ^ cdx_243m ^ cdx_165m ^ cdx_229m ^ cdx_175m ^ cdx_185m ^ cdx_195m ^ cdx_231m ^ cdx_201m ^ r16m;
	reg_0_29 <= cdx_16m ^ cdx_233m ^ cdx_28m ^ cdx_203m ^ cdx_205m ^ cdx_34m ^ cdx_36m ^ cdx_207m ^ cdx_44m ^ cdx_46m ^ cdx_48m ^ cdx_245m ^ cdx_211m ^ cdx_213m ^ cdx_239m ^ cdx_74m ^ cdx_80m ^ cdx_247m ^ cdx_215m ^ cdx_86m ^ cdx_94m ^ cdx_219m ^ cdx_112m ^ cdx_221m ^ cdx_223m ^ cdx_241m ^ cdx_225m ^ cdx_146m ^ cdx_227m ^ cdx_175m ^ cdx_195m ^ cdx_197m ^ cdx_199m ^ r17m;
	reg_0_30 <= cdx_249m ^ cdx_251m ^ cdx_253m ^ cdx_255m ^ cdx_257m ^ cdx_259m ^ cdx_261m ^ cdx_263m ^ cdx_265m ^ cdx_267m ^ cdx_269m ^ cdx_271m ^ cdx_273m ^ cdx_275m ^ cdx_277m ^ cdx_279m ^ cdx_281m ^ cdx_283m ^ cdx_285m ^ cdx_287m ^ cdx_289m ^ cdx_291m ^ cdx_293m ^ cdx_295m ^ cdx_297m ^ cdx_299m ^ cdx_301m ^ cdx_303m ^ cdx_305m ^ r18m;
	reg_0_31 <= cdx_249m ^ cdx_307m ^ cdx_309m ^ cdx_257m ^ cdx_261m ^ cdx_311m ^ cdx_313m ^ cdx_267m ^ cdx_315m ^ cdx_269m ^ cdx_317m ^ cdx_271m ^ cdx_275m ^ cdx_319m ^ cdx_277m ^ cdx_321m ^ cdx_283m ^ cdx_323m ^ cdx_287m ^ cdx_325m ^ cdx_327m ^ cdx_329m ^ cdx_291m ^ cdx_331m ^ cdx_293m ^ cdx_333m ^ cdx_297m ^ cdx_299m ^ cdx_301m ^ cdx_335m ^ r19m;
	reg_0_32 <= cdx_249m ^ cdx_251m ^ cdx_337m ^ cdx_255m ^ cdx_339m ^ cdx_309m ^ cdx_259m ^ cdx_261m ^ cdx_263m ^ cdx_313m ^ cdx_267m ^ cdx_315m ^ cdx_269m ^ cdx_341m ^ cdx_343m ^ cdx_271m ^ cdx_275m ^ cdx_319m ^ cdx_277m ^ cdx_279m ^ cdx_321m ^ cdx_283m ^ cdx_285m ^ cdx_325m ^ cdx_289m ^ cdx_345m ^ cdx_329m ^ cdx_291m ^ cdx_347m ^ cdx_293m ^ cdx_333m ^ cdx_295m ^ cdx_297m ^ cdx_299m ^ cdx_335m ^ cdx_305m ^ r20m;
	reg_0_33 <= cdx_249m ^ cdx_337m ^ cdx_253m ^ cdx_307m ^ cdx_309m ^ cdx_257m ^ cdx_259m ^ cdx_311m ^ cdx_263m ^ cdx_265m ^ cdx_267m ^ cdx_349m ^ cdx_315m ^ cdx_317m ^ cdx_343m ^ cdx_273m ^ cdx_275m ^ cdx_351m ^ cdx_319m ^ cdx_277m ^ cdx_281m ^ cdx_323m ^ cdx_287m ^ cdx_325m ^ cdx_327m ^ cdx_345m ^ cdx_329m ^ cdx_291m ^ cdx_331m ^ cdx_295m ^ cdx_299m ^ cdx_301m ^ cdx_303m ^ r21m;





	reg_1_0 <= a1;
	reg_1_1 <= b1;
	reg_1_2 <= c1;
	reg_1_3 <= d1;
	reg_1_4 <= e1;
	reg_1_5 <= f1;
	reg_1_6 <= g1;
	reg_1_7 <= h1;
	reg_1_8 <= cdx_398m;
	reg_1_9 <= cdx_387m;
	reg_1_10 <= cdx_386m;
	reg_1_11 <= cdx_397m;
	reg_1_12 <= cdx_15m;
	reg_1_13 <= cdx_21m;
	reg_1_14 <= cdx_39m;
	reg_1_15 <= cdx_27m;
	reg_1_16 <= cdx_353m;
	reg_1_17 <= cdx_100m;
	reg_1_18 <= cdx_62m;
	reg_1_19 <= cdx_50m;
	reg_1_20 <= cdx_76m;
	reg_1_21 <= cdx_90m;
	reg_1_22 <= cdx_136m;
	reg_1_23 <= cdx_114m;
	reg_1_24 <= cdx_177m;
	reg_1_25 <= cdx_156m;
	reg_1_26 <= cdx_355m ^ cdx_360m ^ cdx_365m ^ cdx_369m ^ cdx_371m ^ cdx_373m ^ cdx_376m ^ cdx_380m ^ cdx_382m ^ cdx_384m ^ cdx_391m ^ cdx_402m ^ cdx_408m ^ cdx_413m ^ cdx_419m ^ cdx_421m ^ cdx_426m ^ cdx_435m ^ cdx_441m ^ cdx_443m ^ cdx_455m ^ cdx_475m ^ cdx_493m ^ cdx_503m ^ cdx_512m ^ cdx_522m ^ cdx_524m ^ cdx_526m ^ cdx_528m ^ r14m;
	reg_1_27 <= cdx_355m ^ cdx_530m ^ cdx_532m ^ cdx_371m ^ cdx_376m ^ cdx_534m ^ cdx_536m ^ cdx_384m ^ cdx_538m ^ cdx_391m ^ cdx_540m ^ cdx_402m ^ cdx_413m ^ cdx_542m ^ cdx_419m ^ cdx_544m ^ cdx_435m ^ cdx_546m ^ cdx_443m ^ cdx_548m ^ cdx_550m ^ cdx_552m ^ cdx_475m ^ cdx_554m ^ cdx_493m ^ cdx_556m ^ cdx_512m ^ cdx_522m ^ cdx_524m ^ cdx_558m ^ r15m;
	reg_1_28 <= cdx_355m ^ cdx_360m ^ cdx_560m ^ cdx_369m ^ cdx_562m ^ cdx_532m ^ cdx_373m ^ cdx_376m ^ cdx_380m ^ cdx_536m ^ cdx_384m ^ cdx_538m ^ cdx_391m ^ cdx_564m ^ cdx_566m ^ cdx_402m ^ cdx_413m ^ cdx_542m ^ cdx_419m ^ cdx_421m ^ cdx_544m ^ cdx_435m ^ cdx_441m ^ cdx_548m ^ cdx_455m ^ cdx_568m ^ cdx_552m ^ cdx_475m ^ cdx_570m ^ cdx_493m ^ cdx_556m ^ cdx_503m ^ cdx_512m ^ cdx_522m ^ cdx_558m ^ cdx_528m ^ r16m;
	reg_1_29 <= cdx_355m ^ cdx_560m ^ cdx_365m ^ cdx_530m ^ cdx_532m ^ cdx_371m ^ cdx_373m ^ cdx_534m ^ cdx_380m ^ cdx_382m ^ cdx_384m ^ cdx_572m ^ cdx_538m ^ cdx_540m ^ cdx_566m ^ cdx_408m ^ cdx_413m ^ cdx_574m ^ cdx_542m ^ cdx_419m ^ cdx_426m ^ cdx_546m ^ cdx_443m ^ cdx_548m ^ cdx_550m ^ cdx_568m ^ cdx_552m ^ cdx_475m ^ cdx_554m ^ cdx_503m ^ cdx_522m ^ cdx_524m ^ cdx_526m ^ r17m;
	reg_1_30 <= cdx_576m ^ cdx_578m ^ cdx_580m ^ cdx_582m ^ cdx_584m ^ cdx_586m ^ cdx_588m ^ cdx_590m ^ cdx_592m ^ cdx_594m ^ cdx_596m ^ cdx_598m ^ cdx_600m ^ cdx_602m ^ cdx_604m ^ cdx_606m ^ cdx_608m ^ cdx_610m ^ cdx_612m ^ cdx_614m ^ cdx_616m ^ cdx_618m ^ cdx_620m ^ cdx_622m ^ cdx_624m ^ cdx_626m ^ cdx_628m ^ cdx_630m ^ cdx_632m ^ r18m;
	reg_1_31 <= cdx_576m ^ cdx_634m ^ cdx_636m ^ cdx_584m ^ cdx_588m ^ cdx_638m ^ cdx_640m ^ cdx_594m ^ cdx_642m ^ cdx_596m ^ cdx_644m ^ cdx_598m ^ cdx_602m ^ cdx_646m ^ cdx_604m ^ cdx_648m ^ cdx_610m ^ cdx_650m ^ cdx_614m ^ cdx_652m ^ cdx_654m ^ cdx_656m ^ cdx_618m ^ cdx_658m ^ cdx_620m ^ cdx_660m ^ cdx_624m ^ cdx_626m ^ cdx_628m ^ cdx_662m ^ r19m;
	reg_1_32 <= cdx_576m ^ cdx_578m ^ cdx_664m ^ cdx_582m ^ cdx_666m ^ cdx_636m ^ cdx_586m ^ cdx_588m ^ cdx_590m ^ cdx_640m ^ cdx_594m ^ cdx_642m ^ cdx_596m ^ cdx_668m ^ cdx_670m ^ cdx_598m ^ cdx_602m ^ cdx_646m ^ cdx_604m ^ cdx_606m ^ cdx_648m ^ cdx_610m ^ cdx_612m ^ cdx_652m ^ cdx_616m ^ cdx_672m ^ cdx_656m ^ cdx_618m ^ cdx_674m ^ cdx_620m ^ cdx_660m ^ cdx_622m ^ cdx_624m ^ cdx_626m ^ cdx_662m ^ cdx_632m ^ r20m;
	reg_1_33 <= cdx_576m ^ cdx_664m ^ cdx_580m ^ cdx_634m ^ cdx_636m ^ cdx_584m ^ cdx_586m ^ cdx_638m ^ cdx_590m ^ cdx_592m ^ cdx_594m ^ cdx_676m ^ cdx_642m ^ cdx_644m ^ cdx_670m ^ cdx_600m ^ cdx_602m ^ cdx_678m ^ cdx_646m ^ cdx_604m ^ cdx_608m ^ cdx_650m ^ cdx_614m ^ cdx_652m ^ cdx_654m ^ cdx_672m ^ cdx_656m ^ cdx_618m ^ cdx_658m ^ cdx_622m ^ cdx_626m ^ cdx_628m ^ cdx_630m ^ r21m;
end

assign x0 = cdx_19m ^ cdx_25m ^ cdx_31m ^ cdx_33m ^ cdx_35m ^ cdx_37m ^ cdx_43m ^ cdx_45m ^ cdx_47m ^ cdx_49m ^ cdx_61m ^ cdx_73m ^ cdx_75m ^ cdx_85m ^ cdx_87m ^ cdx_89m ^ cdx_99m ^ cdx_109m ^ cdx_111m ^ cdx_113m ^ cdx_135m ^ cdx_155m ^ cdx_174m ^ cdx_176m ^ cdx_194m ^ cdx_196m ^ cdx_198m ^ cdx_200m ^ cdx_202m ^ reg_0_26;
assign y0 = cdx_19m ^ cdx_204m ^ cdx_206m ^ cdx_35m ^ cdx_43m ^ cdx_208m ^ cdx_210m ^ cdx_49m ^ cdx_212m ^ cdx_61m ^ cdx_214m ^ cdx_73m ^ cdx_85m ^ cdx_216m ^ cdx_87m ^ cdx_218m ^ cdx_109m ^ cdx_220m ^ cdx_113m ^ cdx_222m ^ cdx_224m ^ cdx_226m ^ cdx_155m ^ cdx_228m ^ cdx_174m ^ cdx_230m ^ cdx_194m ^ cdx_196m ^ cdx_198m ^ cdx_232m ^ reg_0_27;
assign z0 = cdx_19m ^ cdx_25m ^ cdx_234m ^ cdx_33m ^ cdx_236m ^ cdx_206m ^ cdx_37m ^ cdx_43m ^ cdx_45m ^ cdx_210m ^ cdx_49m ^ cdx_212m ^ cdx_61m ^ cdx_238m ^ cdx_240m ^ cdx_73m ^ cdx_85m ^ cdx_216m ^ cdx_87m ^ cdx_89m ^ cdx_218m ^ cdx_109m ^ cdx_111m ^ cdx_222m ^ cdx_135m ^ cdx_242m ^ cdx_226m ^ cdx_155m ^ cdx_244m ^ cdx_174m ^ cdx_230m ^ cdx_176m ^ cdx_194m ^ cdx_196m ^ cdx_232m ^ cdx_202m ^ reg_0_28;
assign t0 = cdx_19m ^ cdx_234m ^ cdx_31m ^ cdx_204m ^ cdx_206m ^ cdx_35m ^ cdx_37m ^ cdx_208m ^ cdx_45m ^ cdx_47m ^ cdx_49m ^ cdx_246m ^ cdx_212m ^ cdx_214m ^ cdx_240m ^ cdx_75m ^ cdx_85m ^ cdx_248m ^ cdx_216m ^ cdx_87m ^ cdx_99m ^ cdx_220m ^ cdx_113m ^ cdx_222m ^ cdx_224m ^ cdx_242m ^ cdx_226m ^ cdx_155m ^ cdx_228m ^ cdx_176m ^ cdx_196m ^ cdx_198m ^ cdx_200m ^ reg_0_29;
assign m0 = cdx_250m ^ cdx_252m ^ cdx_254m ^ cdx_256m ^ cdx_258m ^ cdx_260m ^ cdx_262m ^ cdx_264m ^ cdx_266m ^ cdx_268m ^ cdx_270m ^ cdx_272m ^ cdx_274m ^ cdx_276m ^ cdx_278m ^ cdx_280m ^ cdx_282m ^ cdx_284m ^ cdx_286m ^ cdx_288m ^ cdx_290m ^ cdx_292m ^ cdx_294m ^ cdx_296m ^ cdx_298m ^ cdx_300m ^ cdx_302m ^ cdx_304m ^ cdx_306m ^ reg_0_30;
assign n0 = cdx_250m ^ cdx_308m ^ cdx_310m ^ cdx_258m ^ cdx_262m ^ cdx_312m ^ cdx_314m ^ cdx_268m ^ cdx_316m ^ cdx_270m ^ cdx_318m ^ cdx_272m ^ cdx_276m ^ cdx_320m ^ cdx_278m ^ cdx_322m ^ cdx_284m ^ cdx_324m ^ cdx_288m ^ cdx_326m ^ cdx_328m ^ cdx_330m ^ cdx_292m ^ cdx_332m ^ cdx_294m ^ cdx_334m ^ cdx_298m ^ cdx_300m ^ cdx_302m ^ cdx_336m ^ reg_0_31;
assign p0 = cdx_250m ^ cdx_252m ^ cdx_338m ^ cdx_256m ^ cdx_340m ^ cdx_310m ^ cdx_260m ^ cdx_262m ^ cdx_264m ^ cdx_314m ^ cdx_268m ^ cdx_316m ^ cdx_270m ^ cdx_342m ^ cdx_344m ^ cdx_272m ^ cdx_276m ^ cdx_320m ^ cdx_278m ^ cdx_280m ^ cdx_322m ^ cdx_284m ^ cdx_286m ^ cdx_326m ^ cdx_290m ^ cdx_346m ^ cdx_330m ^ cdx_292m ^ cdx_348m ^ cdx_294m ^ cdx_334m ^ cdx_296m ^ cdx_298m ^ cdx_300m ^ cdx_336m ^ cdx_306m ^ reg_0_32;
assign q0 = cdx_250m ^ cdx_338m ^ cdx_254m ^ cdx_308m ^ cdx_310m ^ cdx_258m ^ cdx_260m ^ cdx_312m ^ cdx_264m ^ cdx_266m ^ cdx_268m ^ cdx_350m ^ cdx_316m ^ cdx_318m ^ cdx_344m ^ cdx_274m ^ cdx_276m ^ cdx_352m ^ cdx_320m ^ cdx_278m ^ cdx_282m ^ cdx_324m ^ cdx_288m ^ cdx_326m ^ cdx_328m ^ cdx_346m ^ cdx_330m ^ cdx_292m ^ cdx_332m ^ cdx_296m ^ cdx_300m ^ cdx_302m ^ cdx_304m ^ reg_0_33;



assign x1 = cdx_358m ^ cdx_363m ^ cdx_368m ^ cdx_370m ^ cdx_372m ^ cdx_374m ^ cdx_379m ^ cdx_381m ^ cdx_383m ^ cdx_385m ^ cdx_396m ^ cdx_407m ^ cdx_409m ^ cdx_418m ^ cdx_420m ^ cdx_422m ^ cdx_431m ^ cdx_440m ^ cdx_442m ^ cdx_444m ^ cdx_465m ^ cdx_484m ^ cdx_502m ^ cdx_504m ^ cdx_521m ^ cdx_523m ^ cdx_525m ^ cdx_527m ^ cdx_529m ^ reg_1_26;
assign y1 = cdx_358m ^ cdx_531m ^ cdx_533m ^ cdx_372m ^ cdx_379m ^ cdx_535m ^ cdx_537m ^ cdx_385m ^ cdx_539m ^ cdx_396m ^ cdx_541m ^ cdx_407m ^ cdx_418m ^ cdx_543m ^ cdx_420m ^ cdx_545m ^ cdx_440m ^ cdx_547m ^ cdx_444m ^ cdx_549m ^ cdx_551m ^ cdx_553m ^ cdx_484m ^ cdx_555m ^ cdx_502m ^ cdx_557m ^ cdx_521m ^ cdx_523m ^ cdx_525m ^ cdx_559m ^ reg_1_27;
assign z1 = cdx_358m ^ cdx_363m ^ cdx_561m ^ cdx_370m ^ cdx_563m ^ cdx_533m ^ cdx_374m ^ cdx_379m ^ cdx_381m ^ cdx_537m ^ cdx_385m ^ cdx_539m ^ cdx_396m ^ cdx_565m ^ cdx_567m ^ cdx_407m ^ cdx_418m ^ cdx_543m ^ cdx_420m ^ cdx_422m ^ cdx_545m ^ cdx_440m ^ cdx_442m ^ cdx_549m ^ cdx_465m ^ cdx_569m ^ cdx_553m ^ cdx_484m ^ cdx_571m ^ cdx_502m ^ cdx_557m ^ cdx_504m ^ cdx_521m ^ cdx_523m ^ cdx_559m ^ cdx_529m ^ reg_1_28;
assign t1 = cdx_358m ^ cdx_561m ^ cdx_368m ^ cdx_531m ^ cdx_533m ^ cdx_372m ^ cdx_374m ^ cdx_535m ^ cdx_381m ^ cdx_383m ^ cdx_385m ^ cdx_573m ^ cdx_539m ^ cdx_541m ^ cdx_567m ^ cdx_409m ^ cdx_418m ^ cdx_575m ^ cdx_543m ^ cdx_420m ^ cdx_431m ^ cdx_547m ^ cdx_444m ^ cdx_549m ^ cdx_551m ^ cdx_569m ^ cdx_553m ^ cdx_484m ^ cdx_555m ^ cdx_504m ^ cdx_523m ^ cdx_525m ^ cdx_527m ^ reg_1_29;
assign m1 = cdx_577m ^ cdx_579m ^ cdx_581m ^ cdx_583m ^ cdx_585m ^ cdx_587m ^ cdx_589m ^ cdx_591m ^ cdx_593m ^ cdx_595m ^ cdx_597m ^ cdx_599m ^ cdx_601m ^ cdx_603m ^ cdx_605m ^ cdx_607m ^ cdx_609m ^ cdx_611m ^ cdx_613m ^ cdx_615m ^ cdx_617m ^ cdx_619m ^ cdx_621m ^ cdx_623m ^ cdx_625m ^ cdx_627m ^ cdx_629m ^ cdx_631m ^ cdx_633m ^ reg_1_30;
assign n1 = cdx_577m ^ cdx_635m ^ cdx_637m ^ cdx_585m ^ cdx_589m ^ cdx_639m ^ cdx_641m ^ cdx_595m ^ cdx_643m ^ cdx_597m ^ cdx_645m ^ cdx_599m ^ cdx_603m ^ cdx_647m ^ cdx_605m ^ cdx_649m ^ cdx_611m ^ cdx_651m ^ cdx_615m ^ cdx_653m ^ cdx_655m ^ cdx_657m ^ cdx_619m ^ cdx_659m ^ cdx_621m ^ cdx_661m ^ cdx_625m ^ cdx_627m ^ cdx_629m ^ cdx_663m ^ reg_1_31;
assign p1 = cdx_577m ^ cdx_579m ^ cdx_665m ^ cdx_583m ^ cdx_667m ^ cdx_637m ^ cdx_587m ^ cdx_589m ^ cdx_591m ^ cdx_641m ^ cdx_595m ^ cdx_643m ^ cdx_597m ^ cdx_669m ^ cdx_671m ^ cdx_599m ^ cdx_603m ^ cdx_647m ^ cdx_605m ^ cdx_607m ^ cdx_649m ^ cdx_611m ^ cdx_613m ^ cdx_653m ^ cdx_617m ^ cdx_673m ^ cdx_657m ^ cdx_619m ^ cdx_675m ^ cdx_621m ^ cdx_661m ^ cdx_623m ^ cdx_625m ^ cdx_627m ^ cdx_663m ^ cdx_633m ^ reg_1_32;
assign q1 = cdx_577m ^ cdx_665m ^ cdx_581m ^ cdx_635m ^ cdx_637m ^ cdx_585m ^ cdx_587m ^ cdx_639m ^ cdx_591m ^ cdx_593m ^ cdx_595m ^ cdx_677m ^ cdx_643m ^ cdx_645m ^ cdx_671m ^ cdx_601m ^ cdx_603m ^ cdx_679m ^ cdx_647m ^ cdx_605m ^ cdx_609m ^ cdx_651m ^ cdx_615m ^ cdx_653m ^ cdx_655m ^ cdx_673m ^ cdx_657m ^ cdx_619m ^ cdx_659m ^ cdx_623m ^ cdx_627m ^ cdx_629m ^ cdx_631m ^ reg_1_33;



assign x0y0z0t0m0n0p0q0 = {q0,p0,n0,m0,t0,z0,y0,x0};
assign x1y1z1t1m1n1p1q1 = {q1,p1,n1,m1,t1,z1,y1,x1};



endmodule

